
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity ram is
	generic
	(
		DATA_WIDTH : natural := 32;		    -- 4 byte one line of memory
		ADDR_WIDTH : natural := 13			    -- 24576 bytes size of memory
	);

	port(
		i_clk    : in  std_logic;
		i_r_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		i_data   : in  std_logic_vector(DATA_WIDTH-1 downto 0);
		i_we     : in  std_logic;
		i_w_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		o_data   : out std_logic_vector(DATA_WIDTH-1 downto 0)
	);
end entity ram;

architecture arch of ram is

	type ram_t is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(DATA_WIDTH-1 downto 0);


-- GENERATED BY BC_MEM_PACKER

-- DATE: Thu May 18 16:01:02 2017

	signal mem : ram_t := (

--			***** COLOR PALLETE *****

		-- fellas
		0 =>	x"000C4CC8",
		1 =>	x"00A8D8FC",
		2 =>	x"00000000",
		3 =>	x"00EC3820",
		4 =>	x"0000A800",
		5 =>	x"00FCFCFC",
		6 =>	x"00747474",
		7 =>	x"00C0C0C0",
--      Link colors
        8 =>    x"00303030",
        9 =>    x"000CCB83",
        10 =>   x"002C98D8",
        11 =>   x"00004B7B",
        12 =>   x"00FFD9D9",
        13 =>   x"00003299",
        14 =>   x"00B1DFF8",
        15 =>   x"00FFFFFF",
        16 =>   x"008E0018",
        17 =>   x"00FF898E",
        18 =>   x"00000000",
        19 =>   x"00006E8A",
        20 =>   x"00002E55",
        21 =>   x"00CBC74D",
        22 =>   x"00E32F47",
        23 =>   x"00173B00",
        24 =>   x"00007A3E",
        25 =>   x"007ED14A",
        26 =>   x"0000311D",
        27 =>   x"0000675B",
        28 =>   x"000AB4B9",
        29 =>   x"00003D00",
        30 =>   x"00008200",
        31 =>   x"003FD65B",
        32 =>   x"00656565",
        33 =>   x"00B9B9B9",
        34 =>   x"00AFAFAF",
-- 		enemie colors
		35 =>	x"00c0c0c0",
		36 => 	x"000038f8",
		37 => 	x"00bc0000",
		38 =>	x"00ff8868",
		39 => 	x"00ffffff",
																															-- map colors

																															40=> x"00000000",
																															41=> x"00bc0000",
																															42=> x"00d8e800",
																															43=> x"00010100",
																															44=> x"00010000",
																															45=> x"0044a0fc",

							46 => x"00523900",
							47 => x"00271900",
							48 => x"00080400",
							49 => x"00010000",
							50 => x"00d8e800",
							51 => x"00000a00",
							52 => x"0000d600",
							53 => x"00020202",
							54 => x"00010101",
							55 => x"00010100",
							56 => x"00030600",
							57 => x"00105ce4",
							58 => x"0044a0fc",
							59 => x"00bc0000",
							60 => x"005800e4",
							61 => x"00020100",
							62 => x"00f85800",
		63 =>	x"003199FF", -- Unused

            --  ADDED SPRITES HERE
          -- RUPEE SPRITE
		64 => x"0202020F",
		65 => x"3C020202",
		66 => x"02020202",
		67 => x"02020202",
		68 => x"02020F0F",
		69 => x"3C3C0202",
		70 => x"02020202",
		71 => x"02020202",
		72 => x"020F0F0F",
		73 => x"3C3C3C02",
		74 => x"02020202",
		75 => x"02020202",
		76 => x"0F3C0F3C",
		77 => x"023C023C",
		78 => x"02020202",
		79 => x"02020202",
		80 => x"0F0F3C3C",
		81 => x"3C023C3C",
		82 => x"02020202",
		83 => x"02020202",
		84 => x"0F0F3C3C",
		85 => x"3C023C3C",
		86 => x"02020202",
		87 => x"02020202",
		88 => x"0F0F3C3C",
		89 => x"3C023C3C",
		90 => x"02020202",
		91 => x"02020202",
		92 => x"0F0F3C3C",
		93 => x"3C023C3C",
		94 => x"02020202",
		95 => x"02020202",
		96 => x"0F0F3C3C",
		97 => x"3C023C3C",
		98 => x"02020202",
		99 => x"02020202",
		100 => x"0F0F3C3C",
		101 => x"3C023C3C",
		102 => x"02020202",
		103 => x"02020202",
		104 => x"0F0F3C3C",
		105 => x"3C023C3C",
		106 => x"02020202",
		107 => x"02020202",
		108 => x"0F3C0F3C",
		109 => x"3C023C3C",
		110 => x"02020202",
		111 => x"02020202",
		112 => x"3C3C3C0F",
		113 => x"023C023C",
		114 => x"02020202",
		115 => x"02020202",
		116 => x"023C3C3C",
		117 => x"3C3C3C02",
		118 => x"02020202",
		119 => x"02020202",
		120 => x"02023C3C",
		121 => x"3C3C0202",
		122 => x"02020202",
		123 => x"02020202",
		124 => x"0202023C",
		125 => x"3C020202",
		126 => x"02020202",
		127 => x"02020202",

          -- BOMB SPRITE
		128 => x"02020202",
		129 => x"020F0202",
		130 => x"02020202",
		131 => x"02020202",
		132 => x"02020202",
		133 => x"020F0202",
		134 => x"02020202",
		135 => x"02020202",
		136 => x"02020202",
		137 => x"02020F02",
		138 => x"02020202",
		139 => x"02020202",
		140 => x"02020202",
		141 => x"0202020F",
		142 => x"02020202",
		143 => x"02020202",
		144 => x"02020202",
		145 => x"0202020F",
		146 => x"02020202",
		147 => x"02020202",
		148 => x"02020202",
		149 => x"02020F02",
		150 => x"02020202",
		151 => x"02020202",
		152 => x"02020D0D",
		153 => x"0D0D0202",
		154 => x"02020202",
		155 => x"02020202",
		156 => x"020D2E2E",
		157 => x"0D0D0D02",
		158 => x"02020202",
		159 => x"02020202",
		160 => x"0D2E0F2E",
		161 => x"0D0D0D0D",
		162 => x"02020202",
		163 => x"02020202",
		164 => x"0D2E2E0D",
		165 => x"0D0D0D0D",
		166 => x"02020202",
		167 => x"02020202",
		168 => x"0D0D0D0D",
		169 => x"0D0D0D0D",
		170 => x"02020202",
		171 => x"02020202",
		172 => x"0D0D0D0D",
		173 => x"0D0D0D0D",
		174 => x"02020202",
		175 => x"02020202",
		176 => x"020D0D0D",
		177 => x"0D0D0D02",
		178 => x"02020202",
		179 => x"02020202",
		180 => x"02020D0D",
		181 => x"0D0D0202",
		182 => x"02020202",
		183 => x"02020202",
		184 => x"02020202",
		185 => x"02020202",
		186 => x"02020202",
		187 => x"02020202",
		188 => x"02020202",
		189 => x"02020202",
		190 => x"02020202",
		191 => x"02020202",

--			***** 16x16 IMAGES *****
--			OVERWORLD SPRITES


						--  sprite 0
		255 => x"00000000",		-- colors: 40, 40, 40, 40
		256 => x"00000000",		-- colors: 40, 40, 40, 40
		257 => x"00000000",		-- colors: 40, 40, 40, 40
		258 => x"00000000",		-- colors: 40, 40, 40, 40
		259 => x"29292929",		-- colors: 41, 41, 41, 41
		260 => x"29292929",		-- colors: 41, 41, 41, 41
		261 => x"29292929",		-- colors: 41, 41, 41, 41
		262 => x"29292929",		-- colors: 41, 41, 41, 41
		263 => x"00002A2A",		-- colors: 40, 40, 42, 42
		264 => x"2A2A0000",		-- colors: 42, 42, 40, 40
		265 => x"00002A2A",		-- colors: 40, 40, 42, 42
		266 => x"2A2A0000",		-- colors: 42, 42, 40, 40
		267 => x"002A2A2A",		-- colors: 40, 42, 42, 42
		268 => x"2A2A2A00",		-- colors: 42, 42, 42, 40
		269 => x"002A2A2A",		-- colors: 40, 42, 42, 42
		270 => x"2A2A2A00",		-- colors: 42, 42, 42, 40
		271 => x"002A2A2A",		-- colors: 40, 42, 42, 42
		272 => x"2A2A2A00",		-- colors: 42, 42, 42, 40
		273 => x"002A2A2A",		-- colors: 40, 42, 42, 42
		274 => x"2A2A2A00",		-- colors: 42, 42, 42, 40
		275 => x"00002A2A",		-- colors: 40, 40, 42, 42
		276 => x"2A2A0000",		-- colors: 42, 42, 40, 40
		277 => x"00002A2A",		-- colors: 40, 40, 42, 42
		278 => x"2A2A0000",		-- colors: 42, 42, 40, 40
		279 => x"00000000",		-- colors: 40, 40, 40, 40
		280 => x"00000000",		-- colors: 40, 40, 40, 40
		281 => x"00000000",		-- colors: 40, 40, 40, 40
		282 => x"00000000",		-- colors: 40, 40, 40, 40
		283 => x"29292929",		-- colors: 41, 41, 41, 41
		284 => x"29292929",		-- colors: 41, 41, 41, 41
		285 => x"29292929",		-- colors: 41, 41, 41, 41
		286 => x"29292929",		-- colors: 41, 41, 41, 41
		287 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		288 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		289 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		290 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		291 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		292 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		293 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		294 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		295 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		296 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		297 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		298 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		299 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		300 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		301 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		302 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		303 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		304 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		305 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		306 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		307 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		308 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		309 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		310 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		311 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		312 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		313 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		314 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		315 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		316 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		317 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		318 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42

						--  sprite 1
		319 => x"00000000",		-- colors: 40, 40, 40, 40
		320 => x"00000000",		-- colors: 40, 40, 40, 40
		321 => x"00000000",		-- colors: 40, 40, 40, 40
		322 => x"00000000",		-- colors: 40, 40, 40, 40
		323 => x"00000000",		-- colors: 40, 40, 40, 40
		324 => x"00000000",		-- colors: 40, 40, 40, 40
		325 => x"00000000",		-- colors: 40, 40, 40, 40
		326 => x"00000000",		-- colors: 40, 40, 40, 40
		327 => x"00000000",		-- colors: 40, 40, 40, 40
		328 => x"00000000",		-- colors: 40, 40, 40, 40
		329 => x"00000000",		-- colors: 40, 40, 40, 40
		330 => x"00000000",		-- colors: 40, 40, 40, 40
		331 => x"00000000",		-- colors: 40, 40, 40, 40
		332 => x"00000000",		-- colors: 40, 40, 40, 40
		333 => x"00000000",		-- colors: 40, 40, 40, 40
		334 => x"00000000",		-- colors: 40, 40, 40, 40
		335 => x"00000000",		-- colors: 40, 40, 40, 40
		336 => x"00000000",		-- colors: 40, 40, 40, 40
		337 => x"00000000",		-- colors: 40, 40, 40, 40
		338 => x"00000000",		-- colors: 40, 40, 40, 40
		339 => x"00000000",		-- colors: 40, 40, 40, 40
		340 => x"00000000",		-- colors: 40, 40, 40, 40
		341 => x"00000000",		-- colors: 40, 40, 40, 40
		342 => x"00000000",		-- colors: 40, 40, 40, 40
		343 => x"00000000",		-- colors: 40, 40, 40, 40
		344 => x"00000000",		-- colors: 40, 40, 40, 40
		345 => x"00000000",		-- colors: 40, 40, 40, 40
		346 => x"00000000",		-- colors: 40, 40, 40, 40
		347 => x"00000000",		-- colors: 40, 40, 40, 40
		348 => x"00000000",		-- colors: 40, 40, 40, 40
		349 => x"00000000",		-- colors: 40, 40, 40, 40
		350 => x"00000000",		-- colors: 40, 40, 40, 40
		351 => x"29292929",		-- colors: 41, 41, 41, 41
		352 => x"29292929",		-- colors: 41, 41, 41, 41
		353 => x"29292929",		-- colors: 41, 41, 41, 41
		354 => x"29292929",		-- colors: 41, 41, 41, 41
		355 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		356 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		357 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		358 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		359 => x"29290000",		-- colors: 41, 41, 40, 40
		360 => x"00002929",		-- colors: 40, 40, 41, 41
		361 => x"29290000",		-- colors: 41, 41, 40, 40
		362 => x"00002929",		-- colors: 40, 40, 41, 41
		363 => x"29000000",		-- colors: 41, 40, 40, 40
		364 => x"00000029",		-- colors: 40, 40, 40, 41
		365 => x"29000000",		-- colors: 41, 40, 40, 40
		366 => x"00000029",		-- colors: 40, 40, 40, 41
		367 => x"29000000",		-- colors: 41, 40, 40, 40
		368 => x"00000029",		-- colors: 40, 40, 40, 41
		369 => x"29000000",		-- colors: 41, 40, 40, 40
		370 => x"00000029",		-- colors: 40, 40, 40, 41
		371 => x"29290000",		-- colors: 41, 41, 40, 40
		372 => x"00002929",		-- colors: 40, 40, 41, 41
		373 => x"29290000",		-- colors: 41, 41, 40, 40
		374 => x"00002929",		-- colors: 40, 40, 41, 41
		375 => x"29292929",		-- colors: 41, 41, 41, 41
		376 => x"29292929",		-- colors: 41, 41, 41, 41
		377 => x"29292929",		-- colors: 41, 41, 41, 41
		378 => x"29292929",		-- colors: 41, 41, 41, 41
		379 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		380 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		381 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		382 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42

						--  sprite 2
		383 => x"00000000",		-- colors: 40, 40, 40, 40
		384 => x"00000000",		-- colors: 40, 40, 40, 40
		385 => x"29000000",		-- colors: 41, 40, 40, 40
		386 => x"00000029",		-- colors: 40, 40, 40, 41
		387 => x"00000000",		-- colors: 40, 40, 40, 40
		388 => x"00000000",		-- colors: 40, 40, 40, 40
		389 => x"29292929",		-- colors: 41, 41, 41, 41
		390 => x"29292929",		-- colors: 41, 41, 41, 41
		391 => x"00000000",		-- colors: 40, 40, 40, 40
		392 => x"00000000",		-- colors: 40, 40, 40, 40
		393 => x"29000000",		-- colors: 41, 40, 40, 40
		394 => x"00000029",		-- colors: 40, 40, 40, 41
		395 => x"00000000",		-- colors: 40, 40, 40, 40
		396 => x"00000000",		-- colors: 40, 40, 40, 40
		397 => x"29000000",		-- colors: 41, 40, 40, 40
		398 => x"00000029",		-- colors: 40, 40, 40, 41
		399 => x"00000000",		-- colors: 40, 40, 40, 40
		400 => x"00000000",		-- colors: 40, 40, 40, 40
		401 => x"29000000",		-- colors: 41, 40, 40, 40
		402 => x"00000029",		-- colors: 40, 40, 40, 41
		403 => x"00000000",		-- colors: 40, 40, 40, 40
		404 => x"00000000",		-- colors: 40, 40, 40, 40
		405 => x"29292929",		-- colors: 41, 41, 41, 41
		406 => x"29292929",		-- colors: 41, 41, 41, 41
		407 => x"00000000",		-- colors: 40, 40, 40, 40
		408 => x"00000000",		-- colors: 40, 40, 40, 40
		409 => x"29000000",		-- colors: 41, 40, 40, 40
		410 => x"00000029",		-- colors: 40, 40, 40, 41
		411 => x"00000000",		-- colors: 40, 40, 40, 40
		412 => x"00000000",		-- colors: 40, 40, 40, 40
		413 => x"29000000",		-- colors: 41, 40, 40, 40
		414 => x"00000029",		-- colors: 40, 40, 40, 41
		415 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		416 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		417 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		418 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		419 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
		420 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
		421 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
		422 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
		423 => x"2A2A0000",		-- colors: 42, 42, 40, 40
		424 => x"00002A2A",		-- colors: 40, 40, 42, 42
		425 => x"2A2A0000",		-- colors: 42, 42, 40, 40
		426 => x"00002A2A",		-- colors: 40, 40, 42, 42
		427 => x"2A000000",		-- colors: 42, 40, 40, 40
		428 => x"0000002A",		-- colors: 40, 40, 40, 42
		429 => x"2A000000",		-- colors: 42, 40, 40, 40
		430 => x"0000002A",		-- colors: 40, 40, 40, 42
		431 => x"2A000000",		-- colors: 42, 40, 40, 40
		432 => x"0000002A",		-- colors: 40, 40, 40, 42
		433 => x"2A000000",		-- colors: 42, 40, 40, 40
		434 => x"0000002A",		-- colors: 40, 40, 40, 42
		435 => x"2A2A0000",		-- colors: 42, 42, 40, 40
		436 => x"00002A2A",		-- colors: 40, 40, 42, 42
		437 => x"2A2A0000",		-- colors: 42, 42, 40, 40
		438 => x"00002A2A",		-- colors: 40, 40, 42, 42
		439 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		440 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		441 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		442 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		443 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
		444 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
		445 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
		446 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43

						--  sprite 3
		447 => x"00292929",		-- colors: 40, 41, 41, 41
		448 => x"29292900",		-- colors: 41, 41, 41, 40
		449 => x"29292929",		-- colors: 41, 41, 41, 41
		450 => x"29292929",		-- colors: 41, 41, 41, 41
		451 => x"00000000",		-- colors: 40, 40, 40, 40
		452 => x"00000000",		-- colors: 40, 40, 40, 40
		453 => x"29292929",		-- colors: 41, 41, 41, 41
		454 => x"29292929",		-- colors: 41, 41, 41, 41
		455 => x"00292929",		-- colors: 40, 41, 41, 41
		456 => x"29292900",		-- colors: 41, 41, 41, 40
		457 => x"29292929",		-- colors: 41, 41, 41, 41
		458 => x"29292929",		-- colors: 41, 41, 41, 41
		459 => x"00292929",		-- colors: 40, 41, 41, 41
		460 => x"29292900",		-- colors: 41, 41, 41, 40
		461 => x"29292929",		-- colors: 41, 41, 41, 41
		462 => x"29292929",		-- colors: 41, 41, 41, 41
		463 => x"00292929",		-- colors: 40, 41, 41, 41
		464 => x"29292900",		-- colors: 41, 41, 41, 40
		465 => x"29292929",		-- colors: 41, 41, 41, 41
		466 => x"29292929",		-- colors: 41, 41, 41, 41
		467 => x"00000000",		-- colors: 40, 40, 40, 40
		468 => x"00000000",		-- colors: 40, 40, 40, 40
		469 => x"29292929",		-- colors: 41, 41, 41, 41
		470 => x"29292929",		-- colors: 41, 41, 41, 41
		471 => x"00292929",		-- colors: 40, 41, 41, 41
		472 => x"29292900",		-- colors: 41, 41, 41, 40
		473 => x"29292929",		-- colors: 41, 41, 41, 41
		474 => x"29292929",		-- colors: 41, 41, 41, 41
		475 => x"00292929",		-- colors: 40, 41, 41, 41
		476 => x"29292900",		-- colors: 41, 41, 41, 40
		477 => x"29292929",		-- colors: 41, 41, 41, 41
		478 => x"29292929",		-- colors: 41, 41, 41, 41
		479 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		480 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		481 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		482 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		483 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
		484 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
		485 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
		486 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
		487 => x"2A2A2929",		-- colors: 42, 42, 41, 41
		488 => x"29292A2A",		-- colors: 41, 41, 42, 42
		489 => x"2A2A2929",		-- colors: 42, 42, 41, 41
		490 => x"29292A2A",		-- colors: 41, 41, 42, 42
		491 => x"2A292929",		-- colors: 42, 41, 41, 41
		492 => x"2929292A",		-- colors: 41, 41, 41, 42
		493 => x"2A292929",		-- colors: 42, 41, 41, 41
		494 => x"2929292A",		-- colors: 41, 41, 41, 42
		495 => x"2A292929",		-- colors: 42, 41, 41, 41
		496 => x"2929292A",		-- colors: 41, 41, 41, 42
		497 => x"2A292929",		-- colors: 42, 41, 41, 41
		498 => x"2929292A",		-- colors: 41, 41, 41, 42
		499 => x"2A2A2929",		-- colors: 42, 42, 41, 41
		500 => x"29292A2A",		-- colors: 41, 41, 42, 42
		501 => x"2A2A2929",		-- colors: 42, 42, 41, 41
		502 => x"29292A2A",		-- colors: 41, 41, 42, 42
		503 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		504 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		505 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		506 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		507 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
		508 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
		509 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
		510 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43

						--  sprite 4
		511 => x"00292929",		-- colors: 40, 41, 41, 41
		512 => x"29292900",		-- colors: 41, 41, 41, 40
		513 => x"29292929",		-- colors: 41, 41, 41, 41
		514 => x"29292929",		-- colors: 41, 41, 41, 41
		515 => x"00000000",		-- colors: 40, 40, 40, 40
		516 => x"00000000",		-- colors: 40, 40, 40, 40
		517 => x"29292929",		-- colors: 41, 41, 41, 41
		518 => x"29292929",		-- colors: 41, 41, 41, 41
		519 => x"00292929",		-- colors: 40, 41, 41, 41
		520 => x"29292900",		-- colors: 41, 41, 41, 40
		521 => x"29292929",		-- colors: 41, 41, 41, 41
		522 => x"29292929",		-- colors: 41, 41, 41, 41
		523 => x"00292929",		-- colors: 40, 41, 41, 41
		524 => x"29292900",		-- colors: 41, 41, 41, 40
		525 => x"29292929",		-- colors: 41, 41, 41, 41
		526 => x"29292929",		-- colors: 41, 41, 41, 41
		527 => x"00292929",		-- colors: 40, 41, 41, 41
		528 => x"29292900",		-- colors: 41, 41, 41, 40
		529 => x"29292929",		-- colors: 41, 41, 41, 41
		530 => x"29292929",		-- colors: 41, 41, 41, 41
		531 => x"00000000",		-- colors: 40, 40, 40, 40
		532 => x"00000000",		-- colors: 40, 40, 40, 40
		533 => x"29292929",		-- colors: 41, 41, 41, 41
		534 => x"29292929",		-- colors: 41, 41, 41, 41
		535 => x"00292929",		-- colors: 40, 41, 41, 41
		536 => x"29292900",		-- colors: 41, 41, 41, 40
		537 => x"29292929",		-- colors: 41, 41, 41, 41
		538 => x"29292929",		-- colors: 41, 41, 41, 41
		539 => x"00292929",		-- colors: 40, 41, 41, 41
		540 => x"29292900",		-- colors: 41, 41, 41, 40
		541 => x"29292929",		-- colors: 41, 41, 41, 41
		542 => x"29292929",		-- colors: 41, 41, 41, 41
		543 => x"00292929",		-- colors: 40, 41, 41, 41
		544 => x"29292900",		-- colors: 41, 41, 41, 40
		545 => x"29292929",		-- colors: 41, 41, 41, 41
		546 => x"29292929",		-- colors: 41, 41, 41, 41
		547 => x"00000000",		-- colors: 40, 40, 40, 40
		548 => x"00000000",		-- colors: 40, 40, 40, 40
		549 => x"29292929",		-- colors: 41, 41, 41, 41
		550 => x"29292929",		-- colors: 41, 41, 41, 41
		551 => x"00292929",		-- colors: 40, 41, 41, 41
		552 => x"29292900",		-- colors: 41, 41, 41, 40
		553 => x"29292929",		-- colors: 41, 41, 41, 41
		554 => x"29292929",		-- colors: 41, 41, 41, 41
		555 => x"00292929",		-- colors: 40, 41, 41, 41
		556 => x"29292900",		-- colors: 41, 41, 41, 40
		557 => x"29292929",		-- colors: 41, 41, 41, 41
		558 => x"29292929",		-- colors: 41, 41, 41, 41
		559 => x"00292929",		-- colors: 40, 41, 41, 41
		560 => x"29292900",		-- colors: 41, 41, 41, 40
		561 => x"29292929",		-- colors: 41, 41, 41, 41
		562 => x"29292929",		-- colors: 41, 41, 41, 41
		563 => x"00000000",		-- colors: 40, 40, 40, 40
		564 => x"00000000",		-- colors: 40, 40, 40, 40
		565 => x"29292929",		-- colors: 41, 41, 41, 41
		566 => x"29292929",		-- colors: 41, 41, 41, 41
		567 => x"00292929",		-- colors: 40, 41, 41, 41
		568 => x"29292900",		-- colors: 41, 41, 41, 40
		569 => x"29292929",		-- colors: 41, 41, 41, 41
		570 => x"29292929",		-- colors: 41, 41, 41, 41
		571 => x"00292929",		-- colors: 40, 41, 41, 41
		572 => x"29292900",		-- colors: 41, 41, 41, 40
		573 => x"29292929",		-- colors: 41, 41, 41, 41
		574 => x"29292929",		-- colors: 41, 41, 41, 41

						--  sprite 5
		575 => x"00000000",		-- colors: 40, 40, 40, 40
		576 => x"00000000",		-- colors: 40, 40, 40, 40
		577 => x"29000000",		-- colors: 41, 40, 40, 40
		578 => x"00000029",		-- colors: 40, 40, 40, 41
		579 => x"00000000",		-- colors: 40, 40, 40, 40
		580 => x"00000000",		-- colors: 40, 40, 40, 40
		581 => x"29292929",		-- colors: 41, 41, 41, 41
		582 => x"29292929",		-- colors: 41, 41, 41, 41
		583 => x"00000000",		-- colors: 40, 40, 40, 40
		584 => x"00000000",		-- colors: 40, 40, 40, 40
		585 => x"29000000",		-- colors: 41, 40, 40, 40
		586 => x"00000029",		-- colors: 40, 40, 40, 41
		587 => x"00000000",		-- colors: 40, 40, 40, 40
		588 => x"00000000",		-- colors: 40, 40, 40, 40
		589 => x"29000000",		-- colors: 41, 40, 40, 40
		590 => x"00000029",		-- colors: 40, 40, 40, 41
		591 => x"00000000",		-- colors: 40, 40, 40, 40
		592 => x"00000000",		-- colors: 40, 40, 40, 40
		593 => x"29000000",		-- colors: 41, 40, 40, 40
		594 => x"00000029",		-- colors: 40, 40, 40, 41
		595 => x"00000000",		-- colors: 40, 40, 40, 40
		596 => x"00000000",		-- colors: 40, 40, 40, 40
		597 => x"29292929",		-- colors: 41, 41, 41, 41
		598 => x"29292929",		-- colors: 41, 41, 41, 41
		599 => x"00000000",		-- colors: 40, 40, 40, 40
		600 => x"00000000",		-- colors: 40, 40, 40, 40
		601 => x"29000000",		-- colors: 41, 40, 40, 40
		602 => x"00000029",		-- colors: 40, 40, 40, 41
		603 => x"00000000",		-- colors: 40, 40, 40, 40
		604 => x"00000000",		-- colors: 40, 40, 40, 40
		605 => x"29000000",		-- colors: 41, 40, 40, 40
		606 => x"00000029",		-- colors: 40, 40, 40, 41
		607 => x"00000000",		-- colors: 40, 40, 40, 40
		608 => x"00000000",		-- colors: 40, 40, 40, 40
		609 => x"29000000",		-- colors: 41, 40, 40, 40
		610 => x"00000029",		-- colors: 40, 40, 40, 41
		611 => x"00000000",		-- colors: 40, 40, 40, 40
		612 => x"00000000",		-- colors: 40, 40, 40, 40
		613 => x"29292929",		-- colors: 41, 41, 41, 41
		614 => x"29292929",		-- colors: 41, 41, 41, 41
		615 => x"00000000",		-- colors: 40, 40, 40, 40
		616 => x"00000000",		-- colors: 40, 40, 40, 40
		617 => x"29000000",		-- colors: 41, 40, 40, 40
		618 => x"00000029",		-- colors: 40, 40, 40, 41
		619 => x"00000000",		-- colors: 40, 40, 40, 40
		620 => x"00000000",		-- colors: 40, 40, 40, 40
		621 => x"29000000",		-- colors: 41, 40, 40, 40
		622 => x"00000029",		-- colors: 40, 40, 40, 41
		623 => x"00000000",		-- colors: 40, 40, 40, 40
		624 => x"00000000",		-- colors: 40, 40, 40, 40
		625 => x"29000000",		-- colors: 41, 40, 40, 40
		626 => x"00000029",		-- colors: 40, 40, 40, 41
		627 => x"00000000",		-- colors: 40, 40, 40, 40
		628 => x"00000000",		-- colors: 40, 40, 40, 40
		629 => x"29292929",		-- colors: 41, 41, 41, 41
		630 => x"29292929",		-- colors: 41, 41, 41, 41
		631 => x"00000000",		-- colors: 40, 40, 40, 40
		632 => x"00000000",		-- colors: 40, 40, 40, 40
		633 => x"29000000",		-- colors: 41, 40, 40, 40
		634 => x"00000029",		-- colors: 40, 40, 40, 41
		635 => x"00000000",		-- colors: 40, 40, 40, 40
		636 => x"00000000",		-- colors: 40, 40, 40, 40
		637 => x"29000000",		-- colors: 41, 40, 40, 40
		638 => x"00000029",		-- colors: 40, 40, 40, 41

						--  sprite 6
		639 => x"00000000",		-- colors: 40, 40, 40, 40
		640 => x"00000000",		-- colors: 40, 40, 40, 40
		641 => x"00000000",		-- colors: 40, 40, 40, 40
		642 => x"00000000",		-- colors: 40, 40, 40, 40
		643 => x"00000000",		-- colors: 40, 40, 40, 40
		644 => x"00000000",		-- colors: 40, 40, 40, 40
		645 => x"00000000",		-- colors: 40, 40, 40, 40
		646 => x"00000000",		-- colors: 40, 40, 40, 40
		647 => x"00000000",		-- colors: 40, 40, 40, 40
		648 => x"00000000",		-- colors: 40, 40, 40, 40
		649 => x"00000000",		-- colors: 40, 40, 40, 40
		650 => x"00000000",		-- colors: 40, 40, 40, 40
		651 => x"00000000",		-- colors: 40, 40, 40, 40
		652 => x"00000000",		-- colors: 40, 40, 40, 40
		653 => x"00000000",		-- colors: 40, 40, 40, 40
		654 => x"00000000",		-- colors: 40, 40, 40, 40
		655 => x"00000000",		-- colors: 40, 40, 40, 40
		656 => x"00000000",		-- colors: 40, 40, 40, 40
		657 => x"00000000",		-- colors: 40, 40, 40, 40
		658 => x"00000000",		-- colors: 40, 40, 40, 40
		659 => x"00000000",		-- colors: 40, 40, 40, 40
		660 => x"00000000",		-- colors: 40, 40, 40, 40
		661 => x"00000000",		-- colors: 40, 40, 40, 40
		662 => x"00000000",		-- colors: 40, 40, 40, 40
		663 => x"00000000",		-- colors: 40, 40, 40, 40
		664 => x"00000000",		-- colors: 40, 40, 40, 40
		665 => x"00000000",		-- colors: 40, 40, 40, 40
		666 => x"00000000",		-- colors: 40, 40, 40, 40
		667 => x"00000000",		-- colors: 40, 40, 40, 40
		668 => x"00000000",		-- colors: 40, 40, 40, 40
		669 => x"00000000",		-- colors: 40, 40, 40, 40
		670 => x"00000000",		-- colors: 40, 40, 40, 40
		671 => x"00000000",		-- colors: 40, 40, 40, 40
		672 => x"00000000",		-- colors: 40, 40, 40, 40
		673 => x"00000000",		-- colors: 40, 40, 40, 40
		674 => x"00000000",		-- colors: 40, 40, 40, 40
		675 => x"00000000",		-- colors: 40, 40, 40, 40
		676 => x"00000000",		-- colors: 40, 40, 40, 40
		677 => x"00000000",		-- colors: 40, 40, 40, 40
		678 => x"00000000",		-- colors: 40, 40, 40, 40
		679 => x"00000000",		-- colors: 40, 40, 40, 40
		680 => x"00000000",		-- colors: 40, 40, 40, 40
		681 => x"00000000",		-- colors: 40, 40, 40, 40
		682 => x"00000000",		-- colors: 40, 40, 40, 40
		683 => x"00000000",		-- colors: 40, 40, 40, 40
		684 => x"00000000",		-- colors: 40, 40, 40, 40
		685 => x"00000000",		-- colors: 40, 40, 40, 40
		686 => x"00000000",		-- colors: 40, 40, 40, 40
		687 => x"00000000",		-- colors: 40, 40, 40, 40
		688 => x"00000000",		-- colors: 40, 40, 40, 40
		689 => x"00000000",		-- colors: 40, 40, 40, 40
		690 => x"00000000",		-- colors: 40, 40, 40, 40
		691 => x"00000000",		-- colors: 40, 40, 40, 40
		692 => x"00000000",		-- colors: 40, 40, 40, 40
		693 => x"00000000",		-- colors: 40, 40, 40, 40
		694 => x"00000000",		-- colors: 40, 40, 40, 40
		695 => x"00000000",		-- colors: 40, 40, 40, 40
		696 => x"00000000",		-- colors: 40, 40, 40, 40
		697 => x"00000000",		-- colors: 40, 40, 40, 40
		698 => x"00000000",		-- colors: 40, 40, 40, 40
		699 => x"00000000",		-- colors: 40, 40, 40, 40
		700 => x"00000000",		-- colors: 40, 40, 40, 40
		701 => x"00000000",		-- colors: 40, 40, 40, 40
		702 => x"00000000",		-- colors: 40, 40, 40, 40

						--  sprite 7
		703 => x"00000000",		-- colors: 40, 40, 40, 40
		704 => x"00000000",		-- colors: 40, 40, 40, 40
		705 => x"00000000",		-- colors: 40, 40, 40, 40
		706 => x"00000000",		-- colors: 40, 40, 40, 40
		707 => x"29292929",		-- colors: 41, 41, 41, 41
		708 => x"29292929",		-- colors: 41, 41, 41, 41
		709 => x"29292929",		-- colors: 41, 41, 41, 41
		710 => x"29292929",		-- colors: 41, 41, 41, 41
		711 => x"00002A2A",		-- colors: 40, 40, 42, 42
		712 => x"2A2A0000",		-- colors: 42, 42, 40, 40
		713 => x"00002A2A",		-- colors: 40, 40, 42, 42
		714 => x"2A2A0000",		-- colors: 42, 42, 40, 40
		715 => x"002A2A2A",		-- colors: 40, 42, 42, 42
		716 => x"2A2A2A00",		-- colors: 42, 42, 42, 40
		717 => x"002A2A2A",		-- colors: 40, 42, 42, 42
		718 => x"2A2A2A00",		-- colors: 42, 42, 42, 40
		719 => x"002A2A2A",		-- colors: 40, 42, 42, 42
		720 => x"2A2A2A00",		-- colors: 42, 42, 42, 40
		721 => x"002A2A2A",		-- colors: 40, 42, 42, 42
		722 => x"2A2A2A00",		-- colors: 42, 42, 42, 40
		723 => x"00002A2A",		-- colors: 40, 40, 42, 42
		724 => x"2A2A0000",		-- colors: 42, 42, 40, 40
		725 => x"00002A2A",		-- colors: 40, 40, 42, 42
		726 => x"2A2A0000",		-- colors: 42, 42, 40, 40
		727 => x"00000000",		-- colors: 40, 40, 40, 40
		728 => x"00000000",		-- colors: 40, 40, 40, 40
		729 => x"00000000",		-- colors: 40, 40, 40, 40
		730 => x"00000000",		-- colors: 40, 40, 40, 40
		731 => x"29292929",		-- colors: 41, 41, 41, 41
		732 => x"29292929",		-- colors: 41, 41, 41, 41
		733 => x"29292929",		-- colors: 41, 41, 41, 41
		734 => x"29292929",		-- colors: 41, 41, 41, 41
		735 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		736 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		737 => x"2B2A2A2A",		-- colors: 43, 42, 42, 42
		738 => x"2A2A2A2B",		-- colors: 42, 42, 42, 43
		739 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		740 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		741 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
		742 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
		743 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		744 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		745 => x"2B2A2A2A",		-- colors: 43, 42, 42, 42
		746 => x"2A2A2A2B",		-- colors: 42, 42, 42, 43
		747 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		748 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		749 => x"2B2A2A2A",		-- colors: 43, 42, 42, 42
		750 => x"2A2A2A2B",		-- colors: 42, 42, 42, 43
		751 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		752 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		753 => x"2B2A2A2A",		-- colors: 43, 42, 42, 42
		754 => x"2A2A2A2B",		-- colors: 42, 42, 42, 43
		755 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		756 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		757 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
		758 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
		759 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		760 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		761 => x"2B2A2A2A",		-- colors: 43, 42, 42, 42
		762 => x"2A2A2A2B",		-- colors: 42, 42, 42, 43
		763 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		764 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		765 => x"2B2A2A2A",		-- colors: 43, 42, 42, 42
		766 => x"2A2A2A2B",		-- colors: 42, 42, 42, 43

						--  sprite 8
		767 => x"00000000",		-- colors: 40, 40, 40, 40
		768 => x"00000000",		-- colors: 40, 40, 40, 40
		769 => x"00000000",		-- colors: 40, 40, 40, 40
		770 => x"00000000",		-- colors: 40, 40, 40, 40
		771 => x"29292929",		-- colors: 41, 41, 41, 41
		772 => x"29292929",		-- colors: 41, 41, 41, 41
		773 => x"29292929",		-- colors: 41, 41, 41, 41
		774 => x"29292929",		-- colors: 41, 41, 41, 41
		775 => x"00002A2A",		-- colors: 40, 40, 42, 42
		776 => x"2A2A0000",		-- colors: 42, 42, 40, 40
		777 => x"00002A2A",		-- colors: 40, 40, 42, 42
		778 => x"2A2A0000",		-- colors: 42, 42, 40, 40
		779 => x"002A2A2A",		-- colors: 40, 42, 42, 42
		780 => x"2A2A2A00",		-- colors: 42, 42, 42, 40
		781 => x"002A2A2A",		-- colors: 40, 42, 42, 42
		782 => x"2A2A2A00",		-- colors: 42, 42, 42, 40
		783 => x"002A2A2A",		-- colors: 40, 42, 42, 42
		784 => x"2A2A2A00",		-- colors: 42, 42, 42, 40
		785 => x"002A2A2A",		-- colors: 40, 42, 42, 42
		786 => x"2A2A2A00",		-- colors: 42, 42, 42, 40
		787 => x"00002A2A",		-- colors: 40, 40, 42, 42
		788 => x"2A2A0000",		-- colors: 42, 42, 40, 40
		789 => x"00002A2A",		-- colors: 40, 40, 42, 42
		790 => x"2A2A0000",		-- colors: 42, 42, 40, 40
		791 => x"00000000",		-- colors: 40, 40, 40, 40
		792 => x"00000000",		-- colors: 40, 40, 40, 40
		793 => x"00000000",		-- colors: 40, 40, 40, 40
		794 => x"00000000",		-- colors: 40, 40, 40, 40
		795 => x"29292929",		-- colors: 41, 41, 41, 41
		796 => x"29292929",		-- colors: 41, 41, 41, 41
		797 => x"29292929",		-- colors: 41, 41, 41, 41
		798 => x"29292929",		-- colors: 41, 41, 41, 41
		799 => x"2B2A2A2A",		-- colors: 43, 42, 42, 42
		800 => x"2A2A2A2B",		-- colors: 42, 42, 42, 43
		801 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		802 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		803 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
		804 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
		805 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		806 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		807 => x"2B2A2A2A",		-- colors: 43, 42, 42, 42
		808 => x"2A2A2A2B",		-- colors: 42, 42, 42, 43
		809 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		810 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		811 => x"2B2A2A2A",		-- colors: 43, 42, 42, 42
		812 => x"2A2A2A2B",		-- colors: 42, 42, 42, 43
		813 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		814 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		815 => x"2B2A2A2A",		-- colors: 43, 42, 42, 42
		816 => x"2A2A2A2B",		-- colors: 42, 42, 42, 43
		817 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		818 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		819 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
		820 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
		821 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		822 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		823 => x"2B2A2A2A",		-- colors: 43, 42, 42, 42
		824 => x"2A2A2A2B",		-- colors: 42, 42, 42, 43
		825 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		826 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		827 => x"2B2A2A2A",		-- colors: 43, 42, 42, 42
		828 => x"2A2A2A2B",		-- colors: 42, 42, 42, 43
		829 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		830 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42

				----------------------------------------------------

others => x"00000000"
	);


begin

	process(i_clk)
	begin
		if rising_edge(i_clk) then
			-- memory write --
			if i_we = '1' then
				mem(to_integer(unsigned(i_w_addr))) <= i_data;
			end if;
			-- memory read --
			o_data <= mem(to_integer(unsigned(i_r_addr)));

		end if;
	end process;

end architecture arch;
