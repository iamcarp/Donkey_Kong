
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity ram is
	generic
	(
		DATA_WIDTH : natural := 32;		    -- 4 byte one line of memory
		ADDR_WIDTH : natural := 13			    -- 24576 bytes size of memory
	);

	port(
		i_clk    : in  std_logic;
		i_r_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		i_data   : in  std_logic_vector(DATA_WIDTH-1 downto 0);
		i_we     : in  std_logic;
		i_w_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		o_data   : out std_logic_vector(DATA_WIDTH-1 downto 0)
	);
end entity ram;

architecture arch of ram is

	type ram_t is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(DATA_WIDTH-1 downto 0);


-- GENERATED BY BC_MEM_PACKER

-- DATE: Thu May 18 16:01:02 2017

	signal mem : ram_t := (

--			***** COLOR PALLETE *****

		-- fellas
		0 =>	x"000C4CC8", 
		1 =>	x"00A8D8FC", 
		2 =>	x"00000000", 
		3 =>	x"00EC3820", 
		4 =>	x"0000A800", 
		5 =>	x"00FCFCFC", 
		6 =>	x"00747474",
		7 =>	x"00C0C0C0",
--      Link colors
        8 =>    x"00303030",
        9 =>    x"000CCB83",
        10 =>   x"002C98D8", 
        11 =>   x"00004B7B",  
        12 =>   x"00FFD9D9", 
        13 =>   x"00003299", 
        14 =>   x"00B1DFF8", 
        15 =>   x"00FFFFFF", 
        16 =>   x"008E0018", 
        17 =>   x"00FF898E", 
        18 =>   x"00000000", 
        19 =>   x"00006E8A", 
        20 =>   x"00002E55", 
        21 =>   x"00CBC74D", 
        22 =>   x"00E32F47", 
        23 =>   x"00173B00", 
        24 =>   x"00007A3E", 
        25 =>   x"007ED14A", 
        26 =>   x"0000311D", 
        27 =>   x"0000675B", 
        28 =>   x"000AB4B9", 
        29 =>   x"00003D00", 
        30 =>   x"00008200", 
        31 =>   x"003FD65B", 
        32 =>   x"00656565", 
        33 =>   x"00B9B9B9",
        34 =>   x"00AFAFAF",
-- 		enemie colors
		35 =>		x"00c0c0c0",
		36 => 	x"000038f8",
		37 => 	x"00bc0000",
		38 =>		x"00ff8868",
		39 => 	x"00ffffff",
		40 =>		x"0044a0ff",
		41 => 	x"0018f8b8",
		42 => 	x"00003050",
		43 => 	x"00007cac",
		44 =>		x"00105ce4",
		45 =>		x"0000b8f8",
		46 =>		x"00f8b8b8",
		47 =>		x"00000000",
		48 =>		x"00888800",
		49 =>		x"00a8e0ff",
		50 =>		x"0098f858",
		51 =>		x"00005800",
		52 =>		x"0044a800",
		53 =>		x"0064584c",
		54 =>		x"007c7c7c",
		55 =>		x"00584000",
		56 =>		x"00d8e800",
		
			--below not fellas
		57 =>	x"008A7F00", -- R: 0 G: 127 B: 138
		58 =>	x"002E9AFF", -- Unused
		59 =>	x"008D7E00", -- Unused
		60 =>	x"003F95E4", -- Unused
		61 =>	x"003598FF", -- Unused
		62 =>	x"003C9AFC", -- Unused
		63 =>	x"003199FF", -- Unused
		64 =>	x"0069885F", -- Unused
		65 =>	x"00658A6C", -- Unused
		66 =>	x"006A895E", -- Unused
		67 =>	x"003997F7", -- Unused
		68 =>	x"003E95E8", -- Unused
		69 =>	x"003299FF", -- Unused
		70 =>	x"003499FF", -- Unused
		71 =>	x"004A91C0", -- Unused
		72 =>	x"00277FFF", -- Unused
		73 =>	x"00584000", -- Unused
		74 =>	x"00C9DDFF", -- Unused
		75 =>	x"000038F8", -- Unused
		76 =>	x"00007CAC", -- Unused
		77 =>	x"0040A4FF", -- Unused
		78 =>	x"00349DEF", -- Unused
		79 =>	x"003092E0", -- Unused
		80 =>	x"00309AEA", -- Unused
		81 =>	x"00000000", -- Unused
		82 =>	x"00000000", -- Unused
		83 =>	x"00000000", -- Unused
		84 =>	x"00000000", -- Unused
		85 =>	x"00000000", -- Unused
		86 =>	x"00000000", -- Unused
		87 =>	x"00000000", -- Unused
		88 =>	x"00000000", -- Unused
		89 =>	x"00000000", -- Unused
		90 =>	x"00000000", -- Unused
		91 =>	x"00000000", -- Unused
		92 =>	x"00000000", -- Unused
		93 =>	x"00000000", -- Unused
		94 =>	x"00000000", -- Unused
		95 =>	x"00000000", -- Unused
		96 =>	x"00000000", -- Unused
		97 =>	x"00000000", -- Unused
		98 =>	x"00000000", -- Unused
		99 =>	x"00000000", -- Unused
		100 =>	x"00000000", -- Unused
		101 =>	x"00000000", -- Unused
		102 =>	x"00000000", -- Unused
		103 =>	x"00000000", -- Unused
		104 =>	x"00000000", -- Unused
		105 =>	x"00000000", -- Unused
		106 =>	x"00000000", -- Unused
		107 =>	x"00000000", -- Unused
		108 =>	x"00000000", -- Unused
		109 =>	x"00000000", -- Unused
		110 =>	x"00000000", -- Unused
		111 =>	x"00000000", -- Unused
		112 =>	x"00000000", -- Unused
		113 =>	x"00000000", -- Unused
		114 =>	x"00000000", -- Unused
		115 =>	x"00000000", -- Unused
		116 =>	x"00000000", -- Unused
		117 =>	x"00000000", -- Unused
		118 =>	x"00000000", -- Unused
		119 =>	x"00000000", -- Unused
		120 =>	x"00000000", -- Unused
		121 =>	x"00000000", -- Unused
		122 =>	x"00000000", -- Unused
		123 =>	x"00000000", -- Unused
		124 =>	x"00000000", -- Unused
		125 =>	x"00000000", -- Unused
		126 =>	x"00000000", -- Unused
		127 =>	x"00000000", -- Unused
		128 =>	x"00000000", -- Unused
		129 =>	x"00000000", -- Unused
		130 =>	x"00000000", -- Unused
		131 =>	x"00000000", -- Unused
		132 =>	x"00000000", -- Unused
		133 =>	x"00000000", -- Unused
		134 =>	x"00000000", -- Unused
		135 =>	x"00000000", -- Unused
		136 =>	x"00000000", -- Unused
		137 =>	x"00000000", -- Unused
		138 =>	x"00000000", -- Unused
		139 =>	x"00000000", -- Unused
		140 =>	x"00000000", -- Unused
		141 =>	x"00000000", -- Unused
		142 =>	x"00000000", -- Unused
		143 =>	x"00000000", -- Unused
		144 =>	x"00000000", -- Unused
		145 =>	x"00000000", -- Unused
		146 =>	x"00000000", -- Unused
		147 =>	x"00000000", -- Unused
		148 =>	x"00000000", -- Unused
		149 =>	x"00000000", -- Unused
		150 =>	x"00000000", -- Unused
		151 =>	x"00000000", -- Unused
		152 =>	x"00000000", -- Unused
		153 =>	x"00000000", -- Unused
		154 =>	x"00000000", -- Unused
		155 =>	x"00000000", -- Unused
		156 =>	x"00000000", -- Unused
		157 =>	x"00000000", -- Unused
		158 =>	x"00000000", -- Unused
		159 =>	x"00000000", -- Unused
		160 =>	x"00000000", -- Unused
		161 =>	x"00000000", -- Unused
		162 =>	x"00000000", -- Unused
		163 =>	x"00000000", -- Unused
		164 =>	x"00000000", -- Unused
		165 =>	x"00000000", -- Unused
		166 =>	x"00000000", -- Unused
		167 =>	x"00000000", -- Unused
		168 =>	x"00000000", -- Unused
		169 =>	x"00000000", -- Unused
		170 =>	x"00000000", -- Unused
		171 =>	x"00000000", -- Unused
		172 =>	x"00000000", -- Unused
		173 =>	x"00000000", -- Unused
		174 =>	x"00000000", -- Unused
		175 =>	x"00000000", -- Unused
		176 =>	x"00000000", -- Unused
		177 =>	x"00000000", -- Unused
		178 =>	x"00000000", -- Unused
		179 =>	x"00000000", -- Unused
		180 =>	x"00000000", -- Unused
		181 =>	x"00000000", -- Unused
		182 =>	x"00000000", -- Unused
		183 =>	x"00000000", -- Unused
		184 =>	x"00000000", -- Unused
		185 =>	x"00000000", -- Unused
		186 =>	x"00000000", -- Unused
		187 =>	x"00000000", -- Unused
		188 =>	x"00000000", -- Unused
		189 =>	x"00000000", -- Unused
		190 =>	x"00000000", -- Unused
		191 =>	x"00000000", -- Unused
		192 =>	x"00000000", -- Unused
		193 =>	x"00000000", -- Unused
		194 =>	x"00000000", -- Unused
		195 =>	x"00000000", -- Unused
		196 =>	x"00000000", -- Unused
		197 =>	x"00000000", -- Unused
		198 =>	x"00000000", -- Unused
		199 =>	x"00000000", -- Unused
		200 =>	x"00000000", -- Unused
		201 =>	x"00000000", -- Unused
		202 =>	x"00000000", -- Unused
		203 =>	x"00000000", -- Unused
		204 =>	x"00000000", -- Unused
		205 =>	x"00000000", -- Unused
		206 =>	x"00000000", -- Unused
		207 =>	x"00000000", -- Unused
		208 =>	x"00000000", -- Unused
		209 =>	x"00000000", -- Unused
		210 =>	x"00000000", -- Unused
		211 =>	x"00000000", -- Unused
		212 =>	x"00000000", -- Unused
		213 =>	x"00000000", -- Unused
		214 =>	x"00000000", -- Unused
		215 =>	x"00000000", -- Unused
		216 =>	x"00000000", -- Unused
		217 =>	x"00000000", -- Unused
		218 =>	x"00000000", -- Unused
		219 =>	x"00000000", -- Unused
		220 =>	x"00000000", -- Unused
		221 =>	x"00000000", -- Unused
		222 =>	x"00000000", -- Unused
		223 =>	x"00000000", -- Unused
		224 =>	x"00000000", -- Unused
		225 =>	x"00000000", -- Unused
		226 =>	x"00000000", -- Unused
		227 =>	x"00000000", -- Unused
		228 =>	x"00000000", -- Unused
		229 =>	x"00000000", -- Unused
		230 =>	x"00000000", -- Unused
		231 =>	x"00000000", -- Unused
		232 =>	x"00000000", -- Unused
		233 =>	x"00000000", -- Unused
		234 =>	x"00000000", -- Unused
		235 =>	x"00000000", -- Unused
		236 =>	x"00000000", -- Unused
		237 =>	x"00000000", -- Unused
		238 =>	x"00000000", -- Unused
		239 =>	x"00000000", -- Unused
		240 =>	x"00000000", -- Unused
		241 =>	x"00000000", -- Unused
		242 =>	x"00000000", -- Unused
		243 =>	x"00000000", -- Unused
		244 =>	x"00000000", -- Unused
		245 =>	x"00000000", -- Unused
		246 =>	x"00000000", -- Unused
		247 =>	x"00000000", -- Unused
		248 =>	x"00000000", -- Unused
		249 =>	x"00000000", -- Unused
		250 =>	x"00000000", -- Unused
		251 =>	x"00000000", -- Unused
		252 =>	x"00000000", -- Unused
		253 =>	x"00000000", -- Unused
		254 =>	x"00000000", -- Unused

--			***** 16x16 IMAGES *****
--			OVERWORLD SPRITES
                --  sprite 0
        255 => x"00000000",
        256 => x"00000000",
        257 => x"00000000",
        258 => x"00000000",
        259 => x"00020202",
        260 => x"02020202",
        261 => x"02020202",
        262 => x"02020200",
        263 => x"00010102",
        264 => x"02020202",
        265 => x"02020202",
        266 => x"02020200",
        267 => x"00010100",
        268 => x"02020202",
        269 => x"02020202",
        270 => x"02020200",
        271 => x"00010100",
        272 => x"01010102",
        273 => x"02020202",
        274 => x"02020200",
        275 => x"00010100",
        276 => x"01010100",
        277 => x"02020202",
        278 => x"02020200",
        279 => x"00010100",
        280 => x"01010100",
        281 => x"01010102",
        282 => x"02020200",
        283 => x"00010100",
        284 => x"01010100",
        285 => x"01010100",
        286 => x"02020200",
        287 => x"00010100",
        288 => x"01010100",
        289 => x"01010100",
        290 => x"01010100",
        291 => x"00010100",
        292 => x"01010100",
        293 => x"01010100",
        294 => x"01010100",
        295 => x"00010100",
        296 => x"01010100",
        297 => x"01010100",
        298 => x"01010100",
        299 => x"00010100",
        300 => x"01010100",
        301 => x"01010100",
        302 => x"01010100",
        303 => x"00010100",
        304 => x"01010100",
        305 => x"01010100",
        306 => x"01010100",
        307 => x"00010100",
        308 => x"01010100",
        309 => x"01010100",
        310 => x"01010100",
        311 => x"00010100",
        312 => x"01010100",
        313 => x"01010100",
        314 => x"01010100",
        315 => x"00000000",
        316 => x"00000000",
        317 => x"00000000",
        318 => x"00000000",

                --  sprite 1
        319 => x"01010000",
        320 => x"02010101",
        321 => x"01010101",
        322 => x"01010101",
        323 => x"01000000",
        324 => x"00020101",
        325 => x"01010101",
        326 => x"01010101",
        327 => x"01000100",
        328 => x"00020200",
        329 => x"00000202",
        330 => x"01010101",
        331 => x"00010000",
        332 => x"00020100",
        333 => x"00000000",
        334 => x"02010101",
        335 => x"00010000",
        336 => x"00020100",
        337 => x"00000000",
        338 => x"02020101",
        339 => x"00010000",
        340 => x"02010000",
        341 => x"00000000",
        342 => x"00020101",
        343 => x"00000000",
        344 => x"02010000",
        345 => x"02000000",
        346 => x"00020201",
        347 => x"00000000",
        348 => x"02010000",
        349 => x"02000002",
        350 => x"02020201",
        351 => x"01000000",
        352 => x"02010000",
        353 => x"02000002",
        354 => x"00020201",
        355 => x"01000000",
        356 => x"02010000",
        357 => x"02020002",
        358 => x"00020201",
        359 => x"01000000",
        360 => x"02010000",
        361 => x"02020002",
        362 => x"00020201",
        363 => x"00000000",
        364 => x"02000000",
        365 => x"00020002",
        366 => x"02020201",
        367 => x"00000000",
        368 => x"02000000",
        369 => x"00000002",
        370 => x"02000201",
        371 => x"00000000",
        372 => x"00000000",
        373 => x"00020202",
        374 => x"00000101",
        375 => x"01000000",
        376 => x"00000200",
        377 => x"00000202",
        378 => x"02020202",
        379 => x"02020202",
        380 => x"02020202",
        381 => x"02020202",
        382 => x"02020101",

                --  sprite 2
        383 => x"01010101",
        384 => x"01010101",
        385 => x"01010101",
        386 => x"01010101",
        387 => x"01010101",
        388 => x"01010101",
        389 => x"01010101",
        390 => x"01010101",
        391 => x"01010101",
        392 => x"01010101",
        393 => x"01010101",
        394 => x"01010101",
        395 => x"01010101",
        396 => x"01010101",
        397 => x"01010101",
        398 => x"01010101",
        399 => x"01010101",
        400 => x"01010101",
        401 => x"01010101",
        402 => x"01010101",
        403 => x"01010101",
        404 => x"01010101",
        405 => x"01010101",
        406 => x"01010101",
        407 => x"01010101",
        408 => x"01010101",
        409 => x"01010101",
        410 => x"01010101",
        411 => x"01010101",
        412 => x"01010101",
        413 => x"01010101",
        414 => x"01010101",
        415 => x"01010101",
        416 => x"01010101",
        417 => x"01010101",
        418 => x"01010101",
        419 => x"01010101",
        420 => x"01010101",
        421 => x"01010101",
        422 => x"01010101",
        423 => x"01010101",
        424 => x"01010101",
        425 => x"01010101",
        426 => x"01010101",
        427 => x"01010101",
        428 => x"01010101",
        429 => x"01010101",
        430 => x"01010101",
        431 => x"01010101",
        432 => x"01010101",
        433 => x"01010101",
        434 => x"01010101",
        435 => x"01010101",
        436 => x"01010101",
        437 => x"01010101",
        438 => x"01010101",
        439 => x"01010101",
        440 => x"01010101",
        441 => x"01010101",
        442 => x"01010101",
        443 => x"01010101",
        444 => x"01010101",
        445 => x"01010101",
        446 => x"01010101",

                --  sprite 3
        447 => x"01000101",
        448 => x"01030301",
        449 => x"01010100",
        450 => x"01010101",
        451 => x"01000000",
        452 => x"03030303",
        453 => x"01010100",
        454 => x"00020202",
        455 => x"01000000",
        456 => x"00010101",
        457 => x"01010100",
        458 => x"00000002",
        459 => x"01020000",
        460 => x"00010101",
        461 => x"01010100",
        462 => x"02000000",
        463 => x"01030303",
        464 => x"00000001",
        465 => x"01010102",
        466 => x"02000000",
        467 => x"03030303",
        468 => x"03000000",
        469 => x"01010102",
        470 => x"00000000",
        471 => x"01010303",
        472 => x"02000000",
        473 => x"00000102",
        474 => x"00020000",
        475 => x"01010101",
        476 => x"02020000",
        477 => x"00000002",
        478 => x"00020000",
        479 => x"01010101",
        480 => x"01020200",
        481 => x"00000000",
        482 => x"00020000",
        483 => x"01010101",
        484 => x"01010200",
        485 => x"00020000",
        486 => x"02000000",
        487 => x"01010101",
        488 => x"01010202",
        489 => x"00020000",
        490 => x"00020000",
        491 => x"01010101",
        492 => x"01010102",
        493 => x"02020200",
        494 => x"00020000",
        495 => x"01010101",
        496 => x"01010102",
        497 => x"02020202",
        498 => x"00020000",
        499 => x"01010101",
        500 => x"01030303",
        501 => x"03030202",
        502 => x"02020000",
        503 => x"01010101",
        504 => x"03030303",
        505 => x"03030202",
        506 => x"02000000",
        507 => x"01010101",
        508 => x"01010303",
        509 => x"03020202",
        510 => x"02000000",

                --  sprite 4
        511 => x"01020202",
        512 => x"02010101",
        513 => x"01020202",
        514 => x"02020201",
        515 => x"02020202",
        516 => x"02020101",
        517 => x"02020202",
        518 => x"02020202",
        519 => x"02020202",
        520 => x"00020202",
        521 => x"02020202",
        522 => x"02020202",
        523 => x"00020202",
        524 => x"00020202",
        525 => x"02020202",
        526 => x"02020202",
        527 => x"00000000",
        528 => x"00000202",
        529 => x"02020202",
        530 => x"02000000",
        531 => x"00000000",
        532 => x"00000002",
        533 => x"02020200",
        534 => x"00000000",
        535 => x"00000000",
        536 => x"02000000",
        537 => x"02020002",
        538 => x"00000000",
        539 => x"00000000",
        540 => x"02000000",
        541 => x"00000002",
        542 => x"00000002",
        543 => x"00000002",
        544 => x"02020000",
        545 => x"00000202",
        546 => x"02000002",
        547 => x"00000002",
        548 => x"01020000",
        549 => x"00000201",
        550 => x"02000002",
        551 => x"00000002",
        552 => x"01020000",
        553 => x"00000201",
        554 => x"02000002",
        555 => x"00000000",
        556 => x"02000000",
        557 => x"00000002",
        558 => x"00000002",
        559 => x"00000000",
        560 => x"00000000",
        561 => x"00000000",
        562 => x"00000002",
        563 => x"00000002",
        564 => x"02000202",
        565 => x"02020000",
        566 => x"00000002",
        567 => x"00020202",
        568 => x"02000202",
        569 => x"02020202",
        570 => x"00020000",
        571 => x"00020202",
        572 => x"02020202",
        573 => x"02020202",
        574 => x"02020002",

                --  sprite 5
        575 => x"01010101",
        576 => x"01010201",
        577 => x"01010101",
        578 => x"01010101",
        579 => x"01010101",
        580 => x"01020201",
        581 => x"01010101",
        582 => x"01010101",
        583 => x"02020101",
        584 => x"02020201",
        585 => x"01010101",
        586 => x"01010101",
        587 => x"02020202",
        588 => x"02020202",
        589 => x"01010101",
        590 => x"01010101",
        591 => x"02020202",
        592 => x"02020202",
        593 => x"01010101",
        594 => x"01010101",
        595 => x"02020202",
        596 => x"02000202",
        597 => x"01010101",
        598 => x"01010101",
        599 => x"00000202",
        600 => x"00020202",
        601 => x"01010101",
        602 => x"01010101",
        603 => x"00000200",
        604 => x"00020202",
        605 => x"01010101",
        606 => x"01010101",
        607 => x"02000000",
        608 => x"00020202",
        609 => x"01010101",
        610 => x"01010101",
        611 => x"02000000",
        612 => x"02020202",
        613 => x"01010101",
        614 => x"01010101",
        615 => x"00000000",
        616 => x"02020202",
        617 => x"01010101",
        618 => x"01010101",
        619 => x"00000000",
        620 => x"02020200",
        621 => x"01010101",
        622 => x"01010101",
        623 => x"00020000",
        624 => x"00020200",
        625 => x"01010101",
        626 => x"01010101",
        627 => x"00020002",
        628 => x"00020200",
        629 => x"01010101",
        630 => x"01010101",
        631 => x"00020002",
        632 => x"00020200",
        633 => x"01010101",
        634 => x"01010101",
        635 => x"00020000",
        636 => x"02020200",
        637 => x"01010101",
        638 => x"01010101",

                --  sprite 6
        639 => x"01020200",
        640 => x"00000000",
        641 => x"00000000",
        642 => x"00000102",
        643 => x"01020303",
        644 => x"03030303",
        645 => x"03030303",
        646 => x"03030102",
        647 => x"01020303",
        648 => x"03030303",
        649 => x"03030303",
        650 => x"03030102",
        651 => x"01020303",
        652 => x"03030303",
        653 => x"03030303",
        654 => x"03030102",
        655 => x"01020200",
        656 => x"00000000",
        657 => x"00000000",
        658 => x"00000102",
        659 => x"01020303",
        660 => x"03030303",
        661 => x"03030303",
        662 => x"03030102",
        663 => x"01020303",
        664 => x"03030303",
        665 => x"03030303",
        666 => x"03030102",
        667 => x"01020303",
        668 => x"03030303",
        669 => x"03030303",
        670 => x"03030102",
        671 => x"01020200",
        672 => x"00000000",
        673 => x"00000000",
        674 => x"00000102",
        675 => x"01020303",
        676 => x"03030303",
        677 => x"03030303",
        678 => x"03030102",
        679 => x"01020303",
        680 => x"03030303",
        681 => x"03030303",
        682 => x"03030102",
        683 => x"01020303",
        684 => x"03030303",
        685 => x"03030303",
        686 => x"03030102",
        687 => x"01020200",
        688 => x"00000000",
        689 => x"00000000",
        690 => x"00000102",
        691 => x"01020303",
        692 => x"03030303",
        693 => x"03030303",
        694 => x"03030102",
        695 => x"01020303",
        696 => x"03030303",
        697 => x"03030303",
        698 => x"03030102",
        699 => x"01020303",
        700 => x"03030303",
        701 => x"03030303",
        702 => x"03030102",

                --  sprite 7
        703 => x"01010101",
        704 => x"01010101",
        705 => x"01010101",
        706 => x"01010101",
        707 => x"01010101",
        708 => x"00010002",
        709 => x"02020101",
        710 => x"01010101",
        711 => x"01010001",
        712 => x"00000000",
        713 => x"00020202",
        714 => x"02010101",
        715 => x"01010000",
        716 => x"02000000",
        717 => x"00000202",
        718 => x"00020101",
        719 => x"01000000",
        720 => x"00000000",
        721 => x"00000002",
        722 => x"02020101",
        723 => x"01000000",
        724 => x"00000200",
        725 => x"00000200",
        726 => x"02020201",
        727 => x"00000000",
        728 => x"00000000",
        729 => x"00000202",
        730 => x"02020101",
        731 => x"00000200",
        732 => x"00000000",
        733 => x"00000002",
        734 => x"02020201",
        735 => x"01000000",
        736 => x"00000000",
        737 => x"02000002",
        738 => x"02000201",
        739 => x"00000000",
        740 => x"02000000",
        741 => x"00000002",
        742 => x"02020201",
        743 => x"00000000",
        744 => x"00000000",
        745 => x"00020202",
        746 => x"02020101",
        747 => x"00000200",
        748 => x"00000000",
        749 => x"00000200",
        750 => x"02020101",
        751 => x"01000000",
        752 => x"00000002",
        753 => x"02020202",
        754 => x"02010101",
        755 => x"01010100",
        756 => x"00010001",
        757 => x"02020001",
        758 => x"01010101",
        759 => x"01010101",
        760 => x"02010101",
        761 => x"01010202",
        762 => x"02020202",
        763 => x"01010102",
        764 => x"02020202",
        765 => x"02020202",
        766 => x"02020101",

                --  sprite 8
        767 => x"01010002",
        768 => x"01000000",
        769 => x"00010002",
        770 => x"01030101",
        771 => x"01010202",
        772 => x"00000202",
        773 => x"00000202",
        774 => x"01030101",
        775 => x"01010100",
        776 => x"00030202",
        777 => x"03000001",
        778 => x"01030101",
        779 => x"01010100",
        780 => x"00030303",
        781 => x"03000001",
        782 => x"01030101",
        783 => x"00000000",
        784 => x"00000200",
        785 => x"00000002",
        786 => x"01030101",
        787 => x"00020000",
        788 => x"02000202",
        789 => x"02020200",
        790 => x"02030101",
        791 => x"00000000",
        792 => x"00000200",
        793 => x"00000000",
        794 => x"00030201",
        795 => x"00000000",
        796 => x"00000200",
        797 => x"00000002",
        798 => x"00000201",
        799 => x"00000000",
        800 => x"00000200",
        801 => x"00000002",
        802 => x"00000201",
        803 => x"00000000",
        804 => x"00000203",
        805 => x"03000002",
        806 => x"00000201",
        807 => x"00000000",
        808 => x"00000200",
        809 => x"03030303",
        810 => x"02030201",
        811 => x"00000000",
        812 => x"00000203",
        813 => x"03000000",
        814 => x"02030201",
        815 => x"00020000",
        816 => x"02000200",
        817 => x"00000202",
        818 => x"02030201",
        819 => x"00000000",
        820 => x"00000201",
        821 => x"01020000",
        822 => x"00030101",
        823 => x"01020202",
        824 => x"02020202",
        825 => x"02000000",
        826 => x"00030201",
        827 => x"02020202",
        828 => x"02020202",
        829 => x"02020202",
        830 => x"02020202",

                --  sprite 9
        831 => x"01010101",
        832 => x"01010101",
        833 => x"01010202",
        834 => x"00000200",
        835 => x"01010101",
        836 => x"01010101",
        837 => x"01010202",
        838 => x"00000200",
        839 => x"01010101",
        840 => x"01010101",
        841 => x"01010202",
        842 => x"00000200",
        843 => x"01010101",
        844 => x"01010101",
        845 => x"01010002",
        846 => x"00000200",
        847 => x"01010101",
        848 => x"01010101",
        849 => x"01010002",
        850 => x"00000200",
        851 => x"01010101",
        852 => x"01010101",
        853 => x"01010002",
        854 => x"00000200",
        855 => x"01010101",
        856 => x"01010101",
        857 => x"01010002",
        858 => x"00000200",
        859 => x"01010101",
        860 => x"01010101",
        861 => x"01010002",
        862 => x"00000200",
        863 => x"01010101",
        864 => x"01010101",
        865 => x"01000002",
        866 => x"00020200",
        867 => x"01010101",
        868 => x"01010101",
        869 => x"01000202",
        870 => x"00020000",
        871 => x"01010101",
        872 => x"01010101",
        873 => x"01000200",
        874 => x"00020000",
        875 => x"01010101",
        876 => x"01010101",
        877 => x"01000200",
        878 => x"00020000",
        879 => x"01010101",
        880 => x"01010101",
        881 => x"01000200",
        882 => x"00000000",
        883 => x"01010101",
        884 => x"01010101",
        885 => x"00000200",
        886 => x"02000000",
        887 => x"01010101",
        888 => x"01010101",
        889 => x"00000000",
        890 => x"02000000",
        891 => x"01010101",
        892 => x"01010101",
        893 => x"00000101",
        894 => x"00000100",

                --  sprite 10
        895 => x"02020202",
        896 => x"02020202",
        897 => x"02020202",
        898 => x"02020202",
        899 => x"02020202",
        900 => x"02020202",
        901 => x"02020202",
        902 => x"02020202",
        903 => x"02020202",
        904 => x"02020202",
        905 => x"02020202",
        906 => x"02020202",
        907 => x"02020202",
        908 => x"02020202",
        909 => x"02020202",
        910 => x"02020202",
        911 => x"02020202",
        912 => x"02020202",
        913 => x"02020202",
        914 => x"02020202",
        915 => x"02020202",
        916 => x"02020202",
        917 => x"02020202",
        918 => x"02020202",
        919 => x"02020202",
        920 => x"02020202",
        921 => x"02020202",
        922 => x"02020202",
        923 => x"02020202",
        924 => x"02020202",
        925 => x"02020202",
        926 => x"02020202",
        927 => x"02020202",
        928 => x"02020202",
        929 => x"02020202",
        930 => x"02020202",
        931 => x"02020202",
        932 => x"02020202",
        933 => x"02020202",
        934 => x"02020202",
        935 => x"02020202",
        936 => x"02020202",
        937 => x"02020202",
        938 => x"02020202",
        939 => x"02020202",
        940 => x"02020202",
        941 => x"02020202",
        942 => x"02020202",
        943 => x"02020202",
        944 => x"02020202",
        945 => x"02020202",
        946 => x"02020202",
        947 => x"02020202",
        948 => x"02020202",
        949 => x"02020202",
        950 => x"02020202",
        951 => x"02020202",
        952 => x"02020202",
        953 => x"02020202",
        954 => x"02020202",
        955 => x"02020202",
        956 => x"02020202",
        957 => x"02020202",
        958 => x"02020202",

                --  sprite 11
        959 => x"00020000",
        960 => x"02020002",
        961 => x"01010101",
        962 => x"01010002",
        963 => x"00020000",
        964 => x"02020002",
        965 => x"01010101",
        966 => x"01000202",
        967 => x"00020200",
        968 => x"02020002",
        969 => x"01010100",
        970 => x"00000201",
        971 => x"00020200",
        972 => x"02020002",
        973 => x"01010002",
        974 => x"00020303",
        975 => x"00020200",
        976 => x"00020202",
        977 => x"01000200",
        978 => x"02030301",
        979 => x"00020200",
        980 => x"00000202",
        981 => x"00000202",
        982 => x"02010101",
        983 => x"00020200",
        984 => x"02000200",
        985 => x"00020002",
        986 => x"01010101",
        987 => x"00020200",
        988 => x"02000200",
        989 => x"02020002",
        990 => x"01010101",
        991 => x"00020000",
        992 => x"02000200",
        993 => x"02000201",
        994 => x"01010101",
        995 => x"00020002",
        996 => x"02000202",
        997 => x"02020201",
        998 => x"01010101",
        999 => x"00020002",
        1000 => x"00000202",
        1001 => x"00020101",
        1002 => x"01010101",
        1003 => x"00000002",
        1004 => x"00020202",
        1005 => x"00020101",
        1006 => x"01010101",
        1007 => x"00000000",
        1008 => x"00000202",
        1009 => x"02020101",
        1010 => x"01010101",
        1011 => x"00020000",
        1012 => x"00020200",
        1013 => x"02020201",
        1014 => x"01010101",
        1015 => x"00000202",
        1016 => x"02020200",
        1017 => x"02020201",
        1018 => x"01010101",
        1019 => x"00000000",
        1020 => x"00020200",
        1021 => x"02000202",
        1022 => x"01010101",

                --  sprite 12
        1023 => x"01010101",
        1024 => x"01010101",
        1025 => x"01010000",
        1026 => x"02020101",
        1027 => x"01010101",
        1028 => x"01010101",
        1029 => x"01000000",
        1030 => x"00020201",
        1031 => x"01010101",
        1032 => x"01010101",
        1033 => x"00000000",
        1034 => x"00000201",
        1035 => x"01010101",
        1036 => x"01010101",
        1037 => x"01000000",
        1038 => x"00000202",
        1039 => x"01010101",
        1040 => x"01010202",
        1041 => x"01000000",
        1042 => x"00000202",
        1043 => x"01010101",
        1044 => x"01010002",
        1045 => x"01000000",
        1046 => x"00020202",
        1047 => x"01010101",
        1048 => x"01000002",
        1049 => x"01000000",
        1050 => x"00000202",
        1051 => x"01010101",
        1052 => x"01000002",
        1053 => x"02000000",
        1054 => x"00000201",
        1055 => x"01010102",
        1056 => x"02000002",
        1057 => x"00000000",
        1058 => x"00000001",
        1059 => x"01010000",
        1060 => x"02000002",
        1061 => x"00000000",
        1062 => x"00000001",
        1063 => x"01000000",
        1064 => x"00000002",
        1065 => x"00000000",
        1066 => x"00000201",
        1067 => x"01000000",
        1068 => x"02000002",
        1069 => x"01000000",
        1070 => x"00000202",
        1071 => x"01000000",
        1072 => x"02000202",
        1073 => x"02000000",
        1074 => x"00000202",
        1075 => x"01000000",
        1076 => x"02000202",
        1077 => x"00000000",
        1078 => x"00000202",
        1079 => x"00000000",
        1080 => x"00000202",
        1081 => x"02000000",
        1082 => x"00020201",
        1083 => x"00000000",
        1084 => x"00000202",
        1085 => x"02000202",
        1086 => x"00000201",

                --  sprite 13
        1087 => x"01010000",
        1088 => x"02020101",
        1089 => x"01010101",
        1090 => x"01010101",
        1091 => x"01000000",
        1092 => x"00020201",
        1093 => x"01010100",
        1094 => x"02010101",
        1095 => x"00000000",
        1096 => x"00000201",
        1097 => x"01010000",
        1098 => x"00020101",
        1099 => x"01000000",
        1100 => x"00000202",
        1101 => x"01000000",
        1102 => x"00000201",
        1103 => x"01000000",
        1104 => x"00000202",
        1105 => x"02000000",
        1106 => x"00000201",
        1107 => x"01000000",
        1108 => x"00020202",
        1109 => x"01000000",
        1110 => x"00000002",
        1111 => x"01000000",
        1112 => x"00000202",
        1113 => x"01000000",
        1114 => x"00000002",
        1115 => x"02000000",
        1116 => x"00000201",
        1117 => x"01000000",
        1118 => x"00000202",
        1119 => x"00000000",
        1120 => x"00000001",
        1121 => x"00000000",
        1122 => x"00000201",
        1123 => x"00000000",
        1124 => x"00000001",
        1125 => x"00000000",
        1126 => x"00020201",
        1127 => x"00000000",
        1128 => x"00000201",
        1129 => x"00000000",
        1130 => x"00020201",
        1131 => x"01000000",
        1132 => x"00000202",
        1133 => x"01000000",
        1134 => x"00000202",
        1135 => x"02000000",
        1136 => x"00000202",
        1137 => x"02000000",
        1138 => x"00000002",
        1139 => x"00000000",
        1140 => x"00000202",
        1141 => x"01010202",
        1142 => x"00000002",
        1143 => x"02000000",
        1144 => x"00020201",
        1145 => x"00000000",
        1146 => x"02000202",
        1147 => x"02000202",
        1148 => x"00000201",
        1149 => x"00000002",
        1150 => x"02000002",

                --  sprite 14
        1151 => x"01010101",
        1152 => x"01010101",
        1153 => x"01010101",
        1154 => x"01010101",
        1155 => x"01010100",
        1156 => x"02010101",
        1157 => x"01010101",
        1158 => x"01010101",
        1159 => x"01010000",
        1160 => x"00020101",
        1161 => x"01010101",
        1162 => x"01010101",
        1163 => x"01000000",
        1164 => x"00000201",
        1165 => x"01010101",
        1166 => x"01010101",
        1167 => x"02000000",
        1168 => x"00000201",
        1169 => x"01010101",
        1170 => x"01010101",
        1171 => x"01000000",
        1172 => x"00000002",
        1173 => x"01010101",
        1174 => x"01010101",
        1175 => x"01000000",
        1176 => x"00000002",
        1177 => x"00010101",
        1178 => x"01010101",
        1179 => x"01000000",
        1180 => x"00000202",
        1181 => x"00000202",
        1182 => x"02010101",
        1183 => x"00000000",
        1184 => x"00000201",
        1185 => x"00020000",
        1186 => x"00020101",
        1187 => x"00000000",
        1188 => x"00020201",
        1189 => x"00000000",
        1190 => x"00020101",
        1191 => x"00000000",
        1192 => x"00020201",
        1193 => x"00000000",
        1194 => x"00000201",
        1195 => x"01000000",
        1196 => x"00000202",
        1197 => x"01000000",
        1198 => x"00000201",
        1199 => x"02000000",
        1200 => x"00000002",
        1201 => x"01000000",
        1202 => x"00000201",
        1203 => x"01010202",
        1204 => x"00000002",
        1205 => x"01000000",
        1206 => x"00020201",
        1207 => x"00000000",
        1208 => x"02000202",
        1209 => x"01020200",
        1210 => x"00020201",
        1211 => x"00000002",
        1212 => x"02000002",
        1213 => x"01020202",
        1214 => x"00020101",

                --  sprite 15
        1215 => x"01010101",
        1216 => x"01010101",
        1217 => x"01010101",
        1218 => x"01010101",
        1219 => x"01010101",
        1220 => x"01010101",
        1221 => x"01010101",
        1222 => x"01010303",
        1223 => x"01010101",
        1224 => x"01010101",
        1225 => x"01010101",
        1226 => x"01030000",
        1227 => x"01010101",
        1228 => x"01010101",
        1229 => x"01010101",
        1230 => x"01030000",
        1231 => x"01010101",
        1232 => x"01010101",
        1233 => x"01010103",
        1234 => x"03000000",
        1235 => x"01010101",
        1236 => x"01010101",
        1237 => x"01010300",
        1238 => x"00000000",
        1239 => x"01010101",
        1240 => x"01010101",
        1241 => x"01010302",
        1242 => x"03000003",
        1243 => x"01010101",
        1244 => x"01010101",
        1245 => x"01010302",
        1246 => x"03000003",
        1247 => x"01010000",
        1248 => x"00000101",
        1249 => x"01010302",
        1250 => x"03000003",
        1251 => x"01000000",
        1252 => x"00000001",
        1253 => x"01010302",
        1254 => x"03000003",
        1255 => x"00000000",
        1256 => x"00000102",
        1257 => x"01010302",
        1258 => x"03000000",
        1259 => x"00000000",
        1260 => x"00000102",
        1261 => x"01010302",
        1262 => x"03000000",
        1263 => x"00000000",
        1264 => x"00000102",
        1265 => x"01010300",
        1266 => x"00000000",
        1267 => x"00000000",
        1268 => x"00010202",
        1269 => x"01010300",
        1270 => x"00000000",
        1271 => x"01000101",
        1272 => x"01020201",
        1273 => x"01030000",
        1274 => x"00000000",
        1275 => x"01010202",
        1276 => x"02020101",
        1277 => x"03000000",
        1278 => x"00000001",

                --  sprite 16
        1279 => x"01010101",
        1280 => x"01030303",
        1281 => x"03030301",
        1282 => x"01010101",
        1283 => x"03030303",
        1284 => x"03030000",
        1285 => x"00000003",
        1286 => x"03030303",
        1287 => x"00000000",
        1288 => x"00020000",
        1289 => x"00000002",
        1290 => x"00000000",
        1291 => x"00000000",
        1292 => x"00000202",
        1293 => x"02020202",
        1294 => x"00000000",
        1295 => x"00030303",
        1296 => x"03030000",
        1297 => x"00000303",
        1298 => x"03030300",
        1299 => x"03000000",
        1300 => x"00000200",
        1301 => x"00030000",
        1302 => x"00000002",
        1303 => x"00000000",
        1304 => x"00000200",
        1305 => x"00030000",
        1306 => x"00000000",
        1307 => x"02020202",
        1308 => x"02020200",
        1309 => x"00030202",
        1310 => x"02020202",
        1311 => x"00000202",
        1312 => x"02000002",
        1313 => x"00030002",
        1314 => x"02020000",
        1315 => x"00000000",
        1316 => x"00000002",
        1317 => x"00030000",
        1318 => x"00000000",
        1319 => x"02020202",
        1320 => x"02020200",
        1321 => x"00000202",
        1322 => x"02020202",
        1323 => x"00000101",
        1324 => x"01010101",
        1325 => x"01010101",
        1326 => x"01010000",
        1327 => x"00010000",
        1328 => x"02020202",
        1329 => x"02020202",
        1330 => x"00000100",
        1331 => x"01020000",
        1332 => x"02020202",
        1333 => x"02020202",
        1334 => x"00000201",
        1335 => x"01020200",
        1336 => x"02020202",
        1337 => x"02020202",
        1338 => x"00020201",
        1339 => x"02020200",
        1340 => x"02020202",
        1341 => x"02020202",
        1342 => x"00020202",

                --  sprite 17
        1343 => x"01010101",
        1344 => x"01010101",
        1345 => x"01010101",
        1346 => x"01010101",
        1347 => x"03030101",
        1348 => x"01010101",
        1349 => x"01010101",
        1350 => x"01010101",
        1351 => x"00020201",
        1352 => x"01010101",
        1353 => x"01010101",
        1354 => x"01010101",
        1355 => x"00000201",
        1356 => x"01010101",
        1357 => x"01010101",
        1358 => x"01010101",
        1359 => x"00000202",
        1360 => x"02010101",
        1361 => x"01010101",
        1362 => x"01010101",
        1363 => x"00000000",
        1364 => x"02020101",
        1365 => x"01010101",
        1366 => x"01010101",
        1367 => x"02000002",
        1368 => x"03020101",
        1369 => x"01010101",
        1370 => x"01010101",
        1371 => x"02000002",
        1372 => x"03020101",
        1373 => x"01010101",
        1374 => x"01010101",
        1375 => x"02000002",
        1376 => x"03020101",
        1377 => x"01010000",
        1378 => x"00000101",
        1379 => x"02000002",
        1380 => x"03020101",
        1381 => x"01000000",
        1382 => x"00000001",
        1383 => x"00000002",
        1384 => x"03020101",
        1385 => x"00000000",
        1386 => x"00000102",
        1387 => x"00000002",
        1388 => x"03020101",
        1389 => x"00000000",
        1390 => x"00000102",
        1391 => x"00000000",
        1392 => x"00020101",
        1393 => x"00000000",
        1394 => x"00000102",
        1395 => x"00000303",
        1396 => x"02020101",
        1397 => x"00000000",
        1398 => x"00010202",
        1399 => x"00030000",
        1400 => x"00020201",
        1401 => x"01000101",
        1402 => x"01020201",
        1403 => x"01030000",
        1404 => x"00020202",
        1405 => x"01010202",
        1406 => x"02020101",

                --  sprite 18
        1407 => x"00000000",
        1408 => x"01000000",
        1409 => x"02020201",
        1410 => x"00000202",
        1411 => x"00000000",
        1412 => x"01000000",
        1413 => x"00000201",
        1414 => x"00000002",
        1415 => x"00000002",
        1416 => x"01000000",
        1417 => x"00000201",
        1418 => x"00000002",
        1419 => x"00000002",
        1420 => x"01000000",
        1421 => x"00000201",
        1422 => x"00000000",
        1423 => x"00000002",
        1424 => x"01000000",
        1425 => x"00000201",
        1426 => x"00000000",
        1427 => x"00000002",
        1428 => x"01000000",
        1429 => x"00000201",
        1430 => x"00000000",
        1431 => x"02000202",
        1432 => x"01000000",
        1433 => x"00000202",
        1434 => x"01000000",
        1435 => x"01020202",
        1436 => x"01000000",
        1437 => x"00000202",
        1438 => x"02010000",
        1439 => x"01010102",
        1440 => x"02000000",
        1441 => x"00000202",
        1442 => x"02010000",
        1443 => x"01010101",
        1444 => x"02000200",
        1445 => x"00020202",
        1446 => x"02010000",
        1447 => x"01010101",
        1448 => x"01020202",
        1449 => x"02020202",
        1450 => x"02010000",
        1451 => x"01010101",
        1452 => x"01010101",
        1453 => x"02020202",
        1454 => x"02010000",
        1455 => x"01010101",
        1456 => x"01010101",
        1457 => x"01010101",
        1458 => x"02010000",
        1459 => x"01010101",
        1460 => x"01010101",
        1461 => x"01010101",
        1462 => x"01020000",
        1463 => x"01010101",
        1464 => x"01010101",
        1465 => x"01010101",
        1466 => x"01020000",
        1467 => x"01010101",
        1468 => x"01010101",
        1469 => x"01010101",
        1470 => x"01010202",

                --  sprite 19
        1471 => x"00000002",
        1472 => x"01020201",
        1473 => x"00000202",
        1474 => x"01020000",
        1475 => x"00000000",
        1476 => x"02020100",
        1477 => x"00000000",
        1478 => x"02020201",
        1479 => x"00000000",
        1480 => x"02020100",
        1481 => x"00000000",
        1482 => x"02020002",
        1483 => x"01000000",
        1484 => x"02020100",
        1485 => x"00000000",
        1486 => x"00020002",
        1487 => x"01000000",
        1488 => x"02010000",
        1489 => x"00000000",
        1490 => x"00020002",
        1491 => x"00000000",
        1492 => x"02010000",
        1493 => x"00000000",
        1494 => x"00000002",
        1495 => x"00000000",
        1496 => x"02010000",
        1497 => x"00000001",
        1498 => x"01020201",
        1499 => x"00000000",
        1500 => x"02010000",
        1501 => x"00000100",
        1502 => x"00000201",
        1503 => x"00000002",
        1504 => x"02010000",
        1505 => x"00000100",
        1506 => x"00000002",
        1507 => x"00000002",
        1508 => x"02010000",
        1509 => x"00000100",
        1510 => x"00000002",
        1511 => x"01000202",
        1512 => x"02010200",
        1513 => x"00020100",
        1514 => x"00000202",
        1515 => x"01000201",
        1516 => x"01010202",
        1517 => x"00020100",
        1518 => x"00000201",
        1519 => x"00020100",
        1520 => x"00000000",
        1521 => x"02020100",
        1522 => x"00000201",
        1523 => x"00020100",
        1524 => x"00000002",
        1525 => x"02020100",
        1526 => x"00000201",
        1527 => x"00010000",
        1528 => x"00000000",
        1529 => x"02020200",
        1530 => x"00020202",
        1531 => x"02010001",
        1532 => x"00000102",
        1533 => x"01020201",
        1534 => x"01020201",

                --  sprite 20
        1535 => x"01000000",
        1536 => x"00000002",
        1537 => x"02020100",
        1538 => x"00020202",
        1539 => x"01000000",
        1540 => x"00000000",
        1541 => x"02020100",
        1542 => x"00000202",
        1543 => x"01000202",
        1544 => x"00000000",
        1545 => x"02020100",
        1546 => x"00000202",
        1547 => x"01010000",
        1548 => x"02000000",
        1549 => x"02020100",
        1550 => x"00000201",
        1551 => x"01000000",
        1552 => x"02000000",
        1553 => x"02020100",
        1554 => x"00000201",
        1555 => x"01000000",
        1556 => x"02000000",
        1557 => x"02020100",
        1558 => x"02020101",
        1559 => x"01000000",
        1560 => x"02000000",
        1561 => x"02020202",
        1562 => x"01010101",
        1563 => x"01000000",
        1564 => x"02000000",
        1565 => x"02020101",
        1566 => x"01010101",
        1567 => x"01000000",
        1568 => x"02000002",
        1569 => x"02010101",
        1570 => x"01010101",
        1571 => x"01000000",
        1572 => x"02000002",
        1573 => x"02010101",
        1574 => x"01010101",
        1575 => x"02010000",
        1576 => x"02000002",
        1577 => x"02010101",
        1578 => x"01010101",
        1579 => x"02010000",
        1580 => x"02000002",
        1581 => x"02010101",
        1582 => x"01010101",
        1583 => x"02010000",
        1584 => x"02000202",
        1585 => x"01010101",
        1586 => x"01010101",
        1587 => x"02010002",
        1588 => x"02020201",
        1589 => x"01010101",
        1590 => x"01010101",
        1591 => x"02020101",
        1592 => x"01010101",
        1593 => x"01010101",
        1594 => x"01010101",
        1595 => x"01010101",
        1596 => x"01010101",
        1597 => x"01010101",
        1598 => x"01010101",

                --  sprite 21
        1599 => x"00000000",
        1600 => x"00000000",
        1601 => x"03000000",
        1602 => x"00000001",
        1603 => x"02020202",
        1604 => x"02020202",
        1605 => x"03000000",
        1606 => x"00000001",
        1607 => x"01000000",
        1608 => x"00000201",
        1609 => x"03020000",
        1610 => x"00000001",
        1611 => x"01000000",
        1612 => x"00000201",
        1613 => x"03030202",
        1614 => x"02020201",
        1615 => x"01010000",
        1616 => x"00020101",
        1617 => x"03000303",
        1618 => x"03030301",
        1619 => x"01010100",
        1620 => x"02010101",
        1621 => x"03020000",
        1622 => x"00000001",
        1623 => x"01010100",
        1624 => x"02010101",
        1625 => x"03020000",
        1626 => x"00000001",
        1627 => x"01000000",
        1628 => x"00020201",
        1629 => x"03030202",
        1630 => x"02020201",
        1631 => x"01030303",
        1632 => x"03030301",
        1633 => x"03020303",
        1634 => x"03030301",
        1635 => x"03000000",
        1636 => x"00000002",
        1637 => x"03020000",
        1638 => x"00000001",
        1639 => x"03000000",
        1640 => x"00000002",
        1641 => x"03020000",
        1642 => x"00000001",
        1643 => x"03000000",
        1644 => x"00000002",
        1645 => x"03030202",
        1646 => x"02020201",
        1647 => x"03000000",
        1648 => x"00000002",
        1649 => x"03000303",
        1650 => x"03030301",
        1651 => x"03000000",
        1652 => x"00000002",
        1653 => x"03000000",
        1654 => x"00000001",
        1655 => x"03000000",
        1656 => x"00000002",
        1657 => x"02000000",
        1658 => x"00000001",
        1659 => x"02020202",
        1660 => x"02020202",
        1661 => x"02020202",
        1662 => x"02020202",

                --  sprite 22
        1663 => x"01010101",
        1664 => x"01010101",
        1665 => x"01010101",
        1666 => x"01010100",
        1667 => x"01010101",
        1668 => x"01010101",
        1669 => x"01010101",
        1670 => x"00010101",
        1671 => x"01010001",
        1672 => x"01010101",
        1673 => x"01010101",
        1674 => x"01010101",
        1675 => x"01010101",
        1676 => x"01010001",
        1677 => x"01010101",
        1678 => x"01010101",
        1679 => x"01010101",
        1680 => x"01010101",
        1681 => x"01000101",
        1682 => x"01010101",
        1683 => x"01000101",
        1684 => x"01010101",
        1685 => x"01010101",
        1686 => x"01000101",
        1687 => x"01010101",
        1688 => x"01010101",
        1689 => x"01010101",
        1690 => x"01010101",
        1691 => x"01010101",
        1692 => x"00010101",
        1693 => x"01010101",
        1694 => x"01010101",
        1695 => x"01010101",
        1696 => x"01010101",
        1697 => x"01010100",
        1698 => x"01010101",
        1699 => x"01010101",
        1700 => x"01010100",
        1701 => x"01010101",
        1702 => x"01010101",
        1703 => x"01010001",
        1704 => x"01010101",
        1705 => x"01010101",
        1706 => x"01010101",
        1707 => x"01010101",
        1708 => x"01010101",
        1709 => x"01010101",
        1710 => x"01010001",
        1711 => x"01010101",
        1712 => x"01010101",
        1713 => x"01010100",
        1714 => x"01010101",
        1715 => x"00010101",
        1716 => x"01010001",
        1717 => x"01010101",
        1718 => x"01010101",
        1719 => x"01010101",
        1720 => x"01010101",
        1721 => x"01010101",
        1722 => x"01010101",
        1723 => x"01010100",
        1724 => x"01010101",
        1725 => x"01000101",
        1726 => x"01010101",

                --  sprite 23
        1727 => x"03000300",
        1728 => x"02000002",
        1729 => x"00000000",
        1730 => x"00000000",
        1731 => x"03000300",
        1732 => x"02000002",
        1733 => x"02020202",
        1734 => x"02020202",
        1735 => x"03000300",
        1736 => x"02020002",
        1737 => x"01000000",
        1738 => x"00000201",
        1739 => x"02020202",
        1740 => x"02030002",
        1741 => x"01000000",
        1742 => x"00000201",
        1743 => x"03030303",
        1744 => x"03000002",
        1745 => x"01010000",
        1746 => x"00020101",
        1747 => x"03000000",
        1748 => x"00020002",
        1749 => x"01010100",
        1750 => x"02010101",
        1751 => x"03000000",
        1752 => x"00020002",
        1753 => x"01010100",
        1754 => x"02010101",
        1755 => x"02020202",
        1756 => x"02030002",
        1757 => x"01000000",
        1758 => x"00020201",
        1759 => x"03030303",
        1760 => x"03000002",
        1761 => x"01030303",
        1762 => x"03030301",
        1763 => x"03000000",
        1764 => x"00020002",
        1765 => x"03000000",
        1766 => x"00000002",
        1767 => x"03000000",
        1768 => x"00020002",
        1769 => x"03000000",
        1770 => x"00000002",
        1771 => x"02020202",
        1772 => x"02030002",
        1773 => x"03000000",
        1774 => x"00000002",
        1775 => x"03030303",
        1776 => x"03000002",
        1777 => x"03000000",
        1778 => x"00000002",
        1779 => x"03000000",
        1780 => x"00000002",
        1781 => x"03000000",
        1782 => x"00000002",
        1783 => x"03000000",
        1784 => x"00000002",
        1785 => x"03000000",
        1786 => x"00000002",
        1787 => x"02020202",
        1788 => x"02020202",
        1789 => x"02020202",
        1790 => x"02020202",

                --  sprite 24
        1791 => x"01010101",
        1792 => x"01010101",
        1793 => x"01020201",
        1794 => x"01020202",
        1795 => x"01010101",
        1796 => x"01010102",
        1797 => x"02020202",
        1798 => x"02020202",
        1799 => x"01010101",
        1800 => x"01020202",
        1801 => x"02030302",
        1802 => x"02020303",
        1803 => x"01010102",
        1804 => x"02020203",
        1805 => x"03030303",
        1806 => x"03030300",
        1807 => x"01010101",
        1808 => x"02030300",
        1809 => x"03030303",
        1810 => x"03030303",
        1811 => x"01010102",
        1812 => x"02030303",
        1813 => x"03030303",
        1814 => x"00030303",
        1815 => x"01010202",
        1816 => x"03030303",
        1817 => x"03030303",
        1818 => x"03030303",
        1819 => x"01010203",
        1820 => x"03030303",
        1821 => x"03030303",
        1822 => x"03030303",
        1823 => x"01010203",
        1824 => x"03000303",
        1825 => x"03030303",
        1826 => x"03030303",
        1827 => x"01020203",
        1828 => x"03030303",
        1829 => x"03030303",
        1830 => x"03030303",
        1831 => x"01020303",
        1832 => x"03030303",
        1833 => x"03030003",
        1834 => x"03030303",
        1835 => x"01030300",
        1836 => x"03030303",
        1837 => x"03030303",
        1838 => x"03030303",
        1839 => x"01030303",
        1840 => x"03030303",
        1841 => x"03030303",
        1842 => x"03030303",
        1843 => x"01030303",
        1844 => x"03030003",
        1845 => x"03030303",
        1846 => x"03030303",
        1847 => x"01030003",
        1848 => x"03030303",
        1849 => x"00030303",
        1850 => x"03030303",
        1851 => x"01030303",
        1852 => x"03030303",
        1853 => x"03030303",
        1854 => x"03030303",

                --  sprite 25
        1855 => x"01020201",
        1856 => x"01020202",
        1857 => x"01020201",
        1858 => x"01020202",
        1859 => x"02020202",
        1860 => x"02020202",
        1861 => x"02020202",
        1862 => x"02020202",
        1863 => x"02030302",
        1864 => x"02020303",
        1865 => x"02030302",
        1866 => x"02020303",
        1867 => x"03030303",
        1868 => x"03030300",
        1869 => x"03030303",
        1870 => x"03030300",
        1871 => x"03030303",
        1872 => x"03030303",
        1873 => x"03030303",
        1874 => x"03030303",
        1875 => x"03030303",
        1876 => x"00030303",
        1877 => x"03030303",
        1878 => x"00030303",
        1879 => x"03030303",
        1880 => x"03030303",
        1881 => x"03030303",
        1882 => x"03030303",
        1883 => x"03030303",
        1884 => x"03030303",
        1885 => x"03030303",
        1886 => x"03030303",
        1887 => x"03030303",
        1888 => x"03030303",
        1889 => x"03030303",
        1890 => x"03030303",
        1891 => x"03030303",
        1892 => x"03030303",
        1893 => x"03030303",
        1894 => x"03030303",
        1895 => x"03030003",
        1896 => x"03030303",
        1897 => x"03030003",
        1898 => x"03030303",
        1899 => x"03030303",
        1900 => x"03030303",
        1901 => x"03030303",
        1902 => x"03030303",
        1903 => x"03030303",
        1904 => x"03030303",
        1905 => x"03030303",
        1906 => x"03030303",
        1907 => x"03030303",
        1908 => x"03030303",
        1909 => x"03030303",
        1910 => x"03030303",
        1911 => x"00030303",
        1912 => x"03030303",
        1913 => x"00030303",
        1914 => x"03030303",
        1915 => x"03030303",
        1916 => x"03030303",
        1917 => x"03030303",
        1918 => x"03030303",

                --  sprite 26
        1919 => x"01020201",
        1920 => x"01020202",
        1921 => x"02010101",
        1922 => x"01010101",
        1923 => x"02020202",
        1924 => x"02020202",
        1925 => x"02020201",
        1926 => x"01010101",
        1927 => x"02030302",
        1928 => x"02020303",
        1929 => x"03020202",
        1930 => x"02020101",
        1931 => x"03030303",
        1932 => x"03030300",
        1933 => x"03030303",
        1934 => x"02010101",
        1935 => x"03030303",
        1936 => x"03030303",
        1937 => x"03030303",
        1938 => x"01010101",
        1939 => x"03030303",
        1940 => x"00030303",
        1941 => x"03030003",
        1942 => x"01010101",
        1943 => x"03030303",
        1944 => x"03030303",
        1945 => x"03030303",
        1946 => x"02020101",
        1947 => x"03030303",
        1948 => x"03030303",
        1949 => x"03030303",
        1950 => x"03030201",
        1951 => x"03030303",
        1952 => x"03030303",
        1953 => x"00030303",
        1954 => x"03030302",
        1955 => x"03030303",
        1956 => x"03030303",
        1957 => x"03030303",
        1958 => x"00030302",
        1959 => x"03030003",
        1960 => x"03030303",
        1961 => x"03030303",
        1962 => x"03030302",
        1963 => x"03030303",
        1964 => x"03030303",
        1965 => x"03030303",
        1966 => x"03030301",
        1967 => x"03030303",
        1968 => x"03030303",
        1969 => x"03030300",
        1970 => x"03030301",
        1971 => x"03030303",
        1972 => x"03030303",
        1973 => x"03030303",
        1974 => x"03030101",
        1975 => x"00030303",
        1976 => x"03030303",
        1977 => x"03030303",
        1978 => x"03030101",
        1979 => x"03030303",
        1980 => x"03030303",
        1981 => x"03030303",
        1982 => x"03030101",

                --  sprite 27
        1983 => x"01010101",
        1984 => x"01010101",
        1985 => x"01020201",
        1986 => x"01020202",
        1987 => x"01010101",
        1988 => x"01010102",
        1989 => x"02020202",
        1990 => x"02020202",
        1991 => x"01010101",
        1992 => x"01020202",
        1993 => x"02010102",
        1994 => x"02020101",
        1995 => x"01010102",
        1996 => x"02020201",
        1997 => x"01010101",
        1998 => x"01010100",
        1999 => x"01010101",
        2000 => x"02010100",
        2001 => x"01010101",
        2002 => x"01010101",
        2003 => x"01010102",
        2004 => x"02010101",
        2005 => x"01010101",
        2006 => x"00010101",
        2007 => x"01010202",
        2008 => x"01010101",
        2009 => x"01010101",
        2010 => x"01010101",
        2011 => x"01010201",
        2012 => x"01010101",
        2013 => x"01010101",
        2014 => x"01010101",
        2015 => x"01010201",
        2016 => x"01000101",
        2017 => x"01010101",
        2018 => x"01010101",
        2019 => x"01020201",
        2020 => x"01010101",
        2021 => x"01010101",
        2022 => x"01010101",
        2023 => x"01020101",
        2024 => x"01010101",
        2025 => x"01010001",
        2026 => x"01010101",
        2027 => x"01010100",
        2028 => x"01010101",
        2029 => x"01010101",
        2030 => x"01010101",
        2031 => x"01010101",
        2032 => x"01010101",
        2033 => x"01010101",
        2034 => x"01010101",
        2035 => x"01010101",
        2036 => x"01010001",
        2037 => x"01010101",
        2038 => x"01010101",
        2039 => x"01010001",
        2040 => x"01010101",
        2041 => x"00010101",
        2042 => x"01010101",
        2043 => x"01010101",
        2044 => x"01010101",
        2045 => x"01010101",
        2046 => x"01010101",

                --  sprite 28
        2047 => x"01020201",
        2048 => x"01020202",
        2049 => x"01020201",
        2050 => x"01020202",
        2051 => x"02020202",
        2052 => x"02020202",
        2053 => x"02020202",
        2054 => x"02020202",
        2055 => x"02010102",
        2056 => x"02020101",
        2057 => x"02010102",
        2058 => x"02020101",
        2059 => x"01010101",
        2060 => x"01010100",
        2061 => x"01010101",
        2062 => x"01010100",
        2063 => x"01010101",
        2064 => x"01010101",
        2065 => x"01010101",
        2066 => x"01010101",
        2067 => x"01010101",
        2068 => x"00010101",
        2069 => x"01010101",
        2070 => x"00010101",
        2071 => x"01010101",
        2072 => x"01010101",
        2073 => x"01010101",
        2074 => x"01010101",
        2075 => x"01010101",
        2076 => x"01010101",
        2077 => x"01010101",
        2078 => x"01010101",
        2079 => x"01010101",
        2080 => x"01010101",
        2081 => x"01010101",
        2082 => x"01010101",
        2083 => x"01010101",
        2084 => x"01010101",
        2085 => x"01010101",
        2086 => x"01010101",
        2087 => x"01010001",
        2088 => x"01010101",
        2089 => x"01010001",
        2090 => x"01010101",
        2091 => x"01010101",
        2092 => x"01010101",
        2093 => x"01010101",
        2094 => x"01010101",
        2095 => x"01010101",
        2096 => x"01010101",
        2097 => x"01010101",
        2098 => x"01010101",
        2099 => x"01010101",
        2100 => x"01010101",
        2101 => x"01010101",
        2102 => x"01010101",
        2103 => x"00010101",
        2104 => x"01010101",
        2105 => x"00010101",
        2106 => x"01010101",
        2107 => x"01010101",
        2108 => x"01010101",
        2109 => x"01010101",
        2110 => x"01010101",

                --  sprite 29
        2111 => x"01020201",
        2112 => x"01020202",
        2113 => x"02010101",
        2114 => x"01010101",
        2115 => x"02020202",
        2116 => x"02020202",
        2117 => x"02020201",
        2118 => x"01010101",
        2119 => x"02010102",
        2120 => x"02020101",
        2121 => x"01020202",
        2122 => x"02020101",
        2123 => x"01010101",
        2124 => x"01010100",
        2125 => x"01010101",
        2126 => x"02010101",
        2127 => x"01010101",
        2128 => x"01010101",
        2129 => x"01010101",
        2130 => x"01010101",
        2131 => x"01010101",
        2132 => x"00010101",
        2133 => x"01010001",
        2134 => x"01010101",
        2135 => x"01010101",
        2136 => x"01010101",
        2137 => x"01010101",
        2138 => x"02020101",
        2139 => x"01010101",
        2140 => x"01010101",
        2141 => x"01010101",
        2142 => x"01010201",
        2143 => x"01010101",
        2144 => x"01010101",
        2145 => x"00010101",
        2146 => x"01010102",
        2147 => x"01010101",
        2148 => x"01010101",
        2149 => x"01010101",
        2150 => x"00010102",
        2151 => x"01010001",
        2152 => x"01010101",
        2153 => x"01010101",
        2154 => x"01010102",
        2155 => x"01010101",
        2156 => x"01010101",
        2157 => x"01010101",
        2158 => x"01010101",
        2159 => x"01010101",
        2160 => x"01010101",
        2161 => x"01010100",
        2162 => x"01010101",
        2163 => x"01010101",
        2164 => x"01010101",
        2165 => x"01010101",
        2166 => x"01010101",
        2167 => x"00010101",
        2168 => x"01010101",
        2169 => x"01010101",
        2170 => x"01010101",
        2171 => x"01010101",
        2172 => x"01010101",
        2173 => x"01010101",
        2174 => x"01010101",

                --  sprite 30
        2175 => x"01010203",
        2176 => x"03000303",
        2177 => x"03030303",
        2178 => x"03030303",
        2179 => x"01020203",
        2180 => x"03030303",
        2181 => x"03030303",
        2182 => x"03030303",
        2183 => x"01020303",
        2184 => x"03030303",
        2185 => x"03030003",
        2186 => x"03030303",
        2187 => x"01030300",
        2188 => x"03030303",
        2189 => x"03030303",
        2190 => x"03030303",
        2191 => x"01030303",
        2192 => x"03030303",
        2193 => x"03030303",
        2194 => x"03030303",
        2195 => x"01030303",
        2196 => x"03030003",
        2197 => x"03030303",
        2198 => x"03030303",
        2199 => x"01030003",
        2200 => x"03030303",
        2201 => x"00030303",
        2202 => x"03030303",
        2203 => x"01030303",
        2204 => x"03030303",
        2205 => x"03030303",
        2206 => x"03030303",
        2207 => x"03030303",
        2208 => x"03030300",
        2209 => x"03030303",
        2210 => x"03030303",
        2211 => x"03000303",
        2212 => x"03030303",
        2213 => x"03030303",
        2214 => x"00030303",
        2215 => x"03030303",
        2216 => x"03030303",
        2217 => x"03030303",
        2218 => x"03030303",
        2219 => x"03030303",
        2220 => x"03030303",
        2221 => x"03030303",
        2222 => x"03030303",
        2223 => x"01030300",
        2224 => x"03030303",
        2225 => x"03030303",
        2226 => x"03030303",
        2227 => x"01030303",
        2228 => x"03030303",
        2229 => x"03030300",
        2230 => x"03030303",
        2231 => x"01030303",
        2232 => x"03030303",
        2233 => x"03030303",
        2234 => x"03030303",
        2235 => x"01030303",
        2236 => x"03030303",
        2237 => x"03030303",
        2238 => x"03030303",

                --  sprite 31
        2239 => x"03030303",
        2240 => x"03030303",
        2241 => x"03030303",
        2242 => x"03030303",
        2243 => x"03030303",
        2244 => x"03030303",
        2245 => x"03030303",
        2246 => x"03030303",
        2247 => x"03030003",
        2248 => x"03030303",
        2249 => x"03030003",
        2250 => x"03030303",
        2251 => x"03030303",
        2252 => x"03030303",
        2253 => x"03030303",
        2254 => x"03030303",
        2255 => x"03030303",
        2256 => x"03030303",
        2257 => x"03030303",
        2258 => x"03030303",
        2259 => x"03030303",
        2260 => x"03030303",
        2261 => x"03030303",
        2262 => x"03030303",
        2263 => x"00030303",
        2264 => x"03030303",
        2265 => x"00030303",
        2266 => x"03030303",
        2267 => x"03030303",
        2268 => x"03030303",
        2269 => x"03030303",
        2270 => x"03030303",
        2271 => x"03030303",
        2272 => x"03030303",
        2273 => x"03030303",
        2274 => x"03030303",
        2275 => x"03030303",
        2276 => x"00030303",
        2277 => x"03030303",
        2278 => x"00030303",
        2279 => x"03030303",
        2280 => x"03030303",
        2281 => x"03030303",
        2282 => x"03030303",
        2283 => x"03030303",
        2284 => x"03030303",
        2285 => x"03030303",
        2286 => x"03030303",
        2287 => x"03030303",
        2288 => x"03030303",
        2289 => x"03030303",
        2290 => x"03030303",
        2291 => x"03030300",
        2292 => x"03030303",
        2293 => x"03030300",
        2294 => x"03030303",
        2295 => x"03030303",
        2296 => x"03030303",
        2297 => x"03030303",
        2298 => x"03030303",
        2299 => x"03030303",
        2300 => x"03030303",
        2301 => x"03030303",
        2302 => x"03030303",

                --  sprite 32
        2303 => x"03030303",
        2304 => x"03030303",
        2305 => x"00030303",
        2306 => x"03030302",
        2307 => x"03030303",
        2308 => x"03030303",
        2309 => x"03030303",
        2310 => x"00030302",
        2311 => x"03030003",
        2312 => x"03030303",
        2313 => x"03030303",
        2314 => x"03030302",
        2315 => x"03030303",
        2316 => x"03030303",
        2317 => x"03030303",
        2318 => x"03030301",
        2319 => x"03030303",
        2320 => x"03030303",
        2321 => x"03030300",
        2322 => x"03030301",
        2323 => x"03030303",
        2324 => x"03030303",
        2325 => x"03030303",
        2326 => x"03030101",
        2327 => x"00030303",
        2328 => x"03030303",
        2329 => x"03030303",
        2330 => x"03030101",
        2331 => x"03030303",
        2332 => x"03030303",
        2333 => x"03030303",
        2334 => x"03030101",
        2335 => x"03030303",
        2336 => x"03030303",
        2337 => x"03030303",
        2338 => x"00030201",
        2339 => x"03030303",
        2340 => x"00030303",
        2341 => x"03030303",
        2342 => x"03030201",
        2343 => x"03030303",
        2344 => x"03030303",
        2345 => x"03030303",
        2346 => x"03030201",
        2347 => x"03030303",
        2348 => x"03030303",
        2349 => x"03030303",
        2350 => x"03030201",
        2351 => x"03030303",
        2352 => x"03030303",
        2353 => x"03030303",
        2354 => x"03030201",
        2355 => x"03030300",
        2356 => x"03030303",
        2357 => x"03030300",
        2358 => x"03030201",
        2359 => x"03030303",
        2360 => x"03030303",
        2361 => x"03030303",
        2362 => x"03030202",
        2363 => x"03030303",
        2364 => x"03030303",
        2365 => x"03030303",
        2366 => x"03030302",

                --  sprite 33
        2367 => x"01010201",
        2368 => x"01000101",
        2369 => x"01010101",
        2370 => x"01010101",
        2371 => x"01020201",
        2372 => x"01010101",
        2373 => x"01010101",
        2374 => x"01010101",
        2375 => x"01020101",
        2376 => x"01010101",
        2377 => x"01010001",
        2378 => x"01010101",
        2379 => x"01010100",
        2380 => x"01010101",
        2381 => x"01010101",
        2382 => x"01010101",
        2383 => x"01010101",
        2384 => x"01010101",
        2385 => x"01010101",
        2386 => x"01010101",
        2387 => x"01010101",
        2388 => x"01010001",
        2389 => x"01010101",
        2390 => x"01010101",
        2391 => x"01010001",
        2392 => x"01010101",
        2393 => x"00010101",
        2394 => x"01010101",
        2395 => x"01010101",
        2396 => x"01010101",
        2397 => x"01010101",
        2398 => x"01010101",
        2399 => x"01010101",
        2400 => x"01010100",
        2401 => x"01010101",
        2402 => x"01010101",
        2403 => x"01000101",
        2404 => x"01010101",
        2405 => x"01010101",
        2406 => x"00010101",
        2407 => x"01010101",
        2408 => x"01010101",
        2409 => x"01010101",
        2410 => x"01010101",
        2411 => x"01010101",
        2412 => x"01010101",
        2413 => x"01010101",
        2414 => x"01010101",
        2415 => x"01010100",
        2416 => x"01010101",
        2417 => x"01010101",
        2418 => x"01010101",
        2419 => x"01010101",
        2420 => x"01010101",
        2421 => x"01010100",
        2422 => x"01010101",
        2423 => x"01010101",
        2424 => x"01010101",
        2425 => x"01010101",
        2426 => x"01010101",
        2427 => x"01010101",
        2428 => x"01010101",
        2429 => x"01010101",
        2430 => x"01010101",

                --  sprite 34
        2431 => x"01010101",
        2432 => x"01010101",
        2433 => x"01010101",
        2434 => x"01010101",
        2435 => x"01010101",
        2436 => x"01010101",
        2437 => x"01010101",
        2438 => x"01010101",
        2439 => x"01010001",
        2440 => x"01010101",
        2441 => x"01010001",
        2442 => x"01010101",
        2443 => x"01010101",
        2444 => x"01010101",
        2445 => x"01010101",
        2446 => x"01010101",
        2447 => x"01010101",
        2448 => x"01010101",
        2449 => x"01010101",
        2450 => x"01010101",
        2451 => x"01010101",
        2452 => x"01010101",
        2453 => x"01010101",
        2454 => x"01010101",
        2455 => x"00010101",
        2456 => x"01010101",
        2457 => x"00010101",
        2458 => x"01010101",
        2459 => x"01010101",
        2460 => x"01010101",
        2461 => x"01010101",
        2462 => x"01010101",
        2463 => x"01010101",
        2464 => x"01010101",
        2465 => x"01010101",
        2466 => x"01010101",
        2467 => x"01010101",
        2468 => x"00010101",
        2469 => x"01010101",
        2470 => x"00010101",
        2471 => x"01010101",
        2472 => x"01010101",
        2473 => x"01010101",
        2474 => x"01010101",
        2475 => x"01010101",
        2476 => x"01010101",
        2477 => x"01010101",
        2478 => x"01010101",
        2479 => x"01010101",
        2480 => x"01010101",
        2481 => x"01010101",
        2482 => x"01010101",
        2483 => x"01010100",
        2484 => x"01010101",
        2485 => x"01010100",
        2486 => x"01010101",
        2487 => x"01010101",
        2488 => x"01010101",
        2489 => x"01010101",
        2490 => x"01010101",
        2491 => x"01010101",
        2492 => x"01010101",
        2493 => x"01010101",
        2494 => x"01010101",

                --  sprite 35
        2495 => x"01010101",
        2496 => x"01010101",
        2497 => x"00010101",
        2498 => x"01010102",
        2499 => x"01010101",
        2500 => x"01010101",
        2501 => x"01010101",
        2502 => x"00010102",
        2503 => x"01010001",
        2504 => x"01010101",
        2505 => x"01010101",
        2506 => x"01010102",
        2507 => x"01010101",
        2508 => x"01010101",
        2509 => x"01010101",
        2510 => x"01010101",
        2511 => x"01010101",
        2512 => x"01010101",
        2513 => x"01010100",
        2514 => x"01010101",
        2515 => x"01010101",
        2516 => x"01010101",
        2517 => x"01010101",
        2518 => x"01010101",
        2519 => x"00010101",
        2520 => x"01010101",
        2521 => x"01010101",
        2522 => x"01010101",
        2523 => x"01010101",
        2524 => x"01010101",
        2525 => x"01010101",
        2526 => x"01010101",
        2527 => x"01010101",
        2528 => x"01010101",
        2529 => x"01010101",
        2530 => x"00010201",
        2531 => x"01010101",
        2532 => x"00010101",
        2533 => x"01010101",
        2534 => x"01010201",
        2535 => x"01010101",
        2536 => x"01010101",
        2537 => x"01010101",
        2538 => x"01010201",
        2539 => x"01010101",
        2540 => x"01010101",
        2541 => x"01010101",
        2542 => x"01010201",
        2543 => x"01010101",
        2544 => x"01010101",
        2545 => x"01010101",
        2546 => x"01010201",
        2547 => x"01010100",
        2548 => x"01010101",
        2549 => x"01010100",
        2550 => x"01010201",
        2551 => x"01010101",
        2552 => x"01010101",
        2553 => x"01010101",
        2554 => x"01010202",
        2555 => x"01010101",
        2556 => x"01010101",
        2557 => x"01010101",
        2558 => x"01010102",

                --  sprite 36
        2559 => x"03030303",
        2560 => x"03030300",
        2561 => x"03030303",
        2562 => x"03030303",
        2563 => x"03000303",
        2564 => x"03030303",
        2565 => x"03030303",
        2566 => x"00030303",
        2567 => x"03030303",
        2568 => x"03030303",
        2569 => x"03030303",
        2570 => x"03030303",
        2571 => x"03030303",
        2572 => x"03030303",
        2573 => x"03030303",
        2574 => x"03030303",
        2575 => x"01030300",
        2576 => x"03030303",
        2577 => x"03030303",
        2578 => x"03030303",
        2579 => x"01030303",
        2580 => x"03030303",
        2581 => x"03030300",
        2582 => x"03030303",
        2583 => x"01030303",
        2584 => x"03030303",
        2585 => x"03030303",
        2586 => x"03030303",
        2587 => x"01030303",
        2588 => x"03030303",
        2589 => x"03030303",
        2590 => x"03030303",
        2591 => x"01030300",
        2592 => x"03030303",
        2593 => x"03030303",
        2594 => x"03030300",
        2595 => x"01010303",
        2596 => x"03030303",
        2597 => x"03030303",
        2598 => x"03030303",
        2599 => x"01010101",
        2600 => x"03030303",
        2601 => x"00030303",
        2602 => x"03030303",
        2603 => x"01010101",
        2604 => x"01030303",
        2605 => x"03030303",
        2606 => x"03030303",
        2607 => x"01010101",
        2608 => x"02030303",
        2609 => x"03030303",
        2610 => x"03030303",
        2611 => x"01010102",
        2612 => x"02030303",
        2613 => x"03030303",
        2614 => x"03030303",
        2615 => x"01010101",
        2616 => x"01010303",
        2617 => x"00030300",
        2618 => x"03010303",
        2619 => x"01010101",
        2620 => x"01010101",
        2621 => x"03030103",
        2622 => x"01010101",

                --  sprite 37
        2623 => x"03030303",
        2624 => x"03030303",
        2625 => x"03030303",
        2626 => x"03030303",
        2627 => x"03030303",
        2628 => x"00030303",
        2629 => x"03030303",
        2630 => x"00030303",
        2631 => x"03030303",
        2632 => x"03030303",
        2633 => x"03030303",
        2634 => x"03030303",
        2635 => x"03030303",
        2636 => x"03030303",
        2637 => x"03030303",
        2638 => x"03030303",
        2639 => x"03030303",
        2640 => x"03030303",
        2641 => x"03030303",
        2642 => x"03030303",
        2643 => x"03030300",
        2644 => x"03030303",
        2645 => x"03030300",
        2646 => x"03030303",
        2647 => x"03030303",
        2648 => x"03030303",
        2649 => x"03030303",
        2650 => x"03030303",
        2651 => x"03030303",
        2652 => x"03030303",
        2653 => x"03030303",
        2654 => x"03030303",
        2655 => x"03030303",
        2656 => x"03030300",
        2657 => x"03030303",
        2658 => x"03030300",
        2659 => x"03030303",
        2660 => x"03030303",
        2661 => x"03030303",
        2662 => x"03030303",
        2663 => x"00030303",
        2664 => x"03030303",
        2665 => x"00030303",
        2666 => x"03030303",
        2667 => x"03030303",
        2668 => x"03030303",
        2669 => x"03030303",
        2670 => x"03030303",
        2671 => x"03030303",
        2672 => x"03030303",
        2673 => x"03030303",
        2674 => x"03030303",
        2675 => x"03030303",
        2676 => x"03030303",
        2677 => x"03030303",
        2678 => x"03030303",
        2679 => x"00030300",
        2680 => x"03010303",
        2681 => x"00030300",
        2682 => x"03010303",
        2683 => x"03030103",
        2684 => x"01010101",
        2685 => x"03030103",
        2686 => x"01010101",

                --  sprite 38
        2687 => x"03030303",
        2688 => x"03030303",
        2689 => x"03030303",
        2690 => x"00030201",
        2691 => x"03030303",
        2692 => x"00030303",
        2693 => x"03030303",
        2694 => x"03030201",
        2695 => x"03030303",
        2696 => x"03030303",
        2697 => x"03030303",
        2698 => x"03030201",
        2699 => x"03030303",
        2700 => x"03030303",
        2701 => x"03030303",
        2702 => x"03030201",
        2703 => x"03030303",
        2704 => x"03030303",
        2705 => x"03030303",
        2706 => x"03030201",
        2707 => x"03030300",
        2708 => x"03030303",
        2709 => x"03030300",
        2710 => x"03030201",
        2711 => x"03030303",
        2712 => x"03030303",
        2713 => x"03030303",
        2714 => x"03030202",
        2715 => x"03030303",
        2716 => x"03030303",
        2717 => x"03030303",
        2718 => x"03030302",
        2719 => x"03030303",
        2720 => x"03030300",
        2721 => x"03030303",
        2722 => x"03030301",
        2723 => x"03030303",
        2724 => x"03030303",
        2725 => x"03000303",
        2726 => x"03000301",
        2727 => x"00030303",
        2728 => x"03030303",
        2729 => x"03030303",
        2730 => x"03030101",
        2731 => x"03030303",
        2732 => x"03030303",
        2733 => x"03030303",
        2734 => x"01010101",
        2735 => x"03030303",
        2736 => x"03030303",
        2737 => x"03030303",
        2738 => x"02010101",
        2739 => x"03030303",
        2740 => x"03030303",
        2741 => x"00030303",
        2742 => x"02020101",
        2743 => x"00030300",
        2744 => x"03010303",
        2745 => x"03030301",
        2746 => x"01010101",
        2747 => x"03030103",
        2748 => x"01010101",
        2749 => x"01010101",
        2750 => x"01010101",

                --  sprite 39
        2751 => x"01010101",
        2752 => x"01010100",
        2753 => x"01010101",
        2754 => x"01010101",
        2755 => x"01000101",
        2756 => x"01010101",
        2757 => x"01010101",
        2758 => x"00010101",
        2759 => x"01010101",
        2760 => x"01010101",
        2761 => x"01010101",
        2762 => x"01010101",
        2763 => x"01010101",
        2764 => x"01010101",
        2765 => x"01010101",
        2766 => x"01010101",
        2767 => x"01010100",
        2768 => x"01010101",
        2769 => x"01010101",
        2770 => x"01010101",
        2771 => x"01010101",
        2772 => x"01010101",
        2773 => x"01010100",
        2774 => x"01010101",
        2775 => x"01010101",
        2776 => x"01010101",
        2777 => x"01010101",
        2778 => x"01010101",
        2779 => x"01010101",
        2780 => x"01010101",
        2781 => x"01010101",
        2782 => x"01010101",
        2783 => x"01010100",
        2784 => x"01010101",
        2785 => x"01010101",
        2786 => x"01010100",
        2787 => x"01010101",
        2788 => x"01010101",
        2789 => x"01010101",
        2790 => x"01010101",
        2791 => x"01010101",
        2792 => x"01010101",
        2793 => x"00010101",
        2794 => x"01010101",
        2795 => x"01010101",
        2796 => x"01010101",
        2797 => x"01010101",
        2798 => x"01010101",
        2799 => x"01010101",
        2800 => x"02010101",
        2801 => x"01010101",
        2802 => x"01010101",
        2803 => x"01010102",
        2804 => x"02010101",
        2805 => x"01010101",
        2806 => x"01010101",
        2807 => x"01010101",
        2808 => x"01010101",
        2809 => x"00010100",
        2810 => x"01010101",
        2811 => x"01010101",
        2812 => x"01010101",
        2813 => x"01010101",
        2814 => x"01010101",

                --  sprite 40
        2815 => x"01010101",
        2816 => x"01010101",
        2817 => x"01010101",
        2818 => x"01010101",
        2819 => x"01010101",
        2820 => x"00010101",
        2821 => x"01010101",
        2822 => x"00010101",
        2823 => x"01010101",
        2824 => x"01010101",
        2825 => x"01010101",
        2826 => x"01010101",
        2827 => x"01010101",
        2828 => x"01010101",
        2829 => x"01010101",
        2830 => x"01010101",
        2831 => x"01010101",
        2832 => x"01010101",
        2833 => x"01010101",
        2834 => x"01010101",
        2835 => x"01010100",
        2836 => x"01010101",
        2837 => x"01010100",
        2838 => x"01010101",
        2839 => x"01010101",
        2840 => x"01010101",
        2841 => x"01010101",
        2842 => x"01010101",
        2843 => x"01010101",
        2844 => x"01010101",
        2845 => x"01010101",
        2846 => x"01010101",
        2847 => x"01010101",
        2848 => x"01010100",
        2849 => x"01010101",
        2850 => x"01010100",
        2851 => x"01010101",
        2852 => x"01010101",
        2853 => x"01010101",
        2854 => x"01010101",
        2855 => x"00010101",
        2856 => x"01010101",
        2857 => x"00010101",
        2858 => x"01010101",
        2859 => x"01010101",
        2860 => x"01010101",
        2861 => x"01010101",
        2862 => x"01010101",
        2863 => x"01010101",
        2864 => x"01010101",
        2865 => x"01010101",
        2866 => x"01010101",
        2867 => x"01010101",
        2868 => x"01010101",
        2869 => x"01010101",
        2870 => x"01010101",
        2871 => x"00010100",
        2872 => x"01010101",
        2873 => x"00010100",
        2874 => x"01010101",
        2875 => x"01010101",
        2876 => x"01010101",
        2877 => x"01010101",
        2878 => x"01010101",

                --  sprite 41
        2879 => x"01010101",
        2880 => x"01010101",
        2881 => x"01010101",
        2882 => x"00010201",
        2883 => x"01010101",
        2884 => x"00010101",
        2885 => x"01010101",
        2886 => x"01010201",
        2887 => x"01010101",
        2888 => x"01010101",
        2889 => x"01010101",
        2890 => x"01010201",
        2891 => x"01010101",
        2892 => x"01010101",
        2893 => x"01010101",
        2894 => x"01010201",
        2895 => x"01010101",
        2896 => x"01010101",
        2897 => x"01010101",
        2898 => x"01010201",
        2899 => x"01010100",
        2900 => x"01010101",
        2901 => x"01010100",
        2902 => x"01010201",
        2903 => x"01010101",
        2904 => x"01010101",
        2905 => x"01010101",
        2906 => x"01010202",
        2907 => x"01010101",
        2908 => x"01010101",
        2909 => x"01010101",
        2910 => x"01010102",
        2911 => x"01010101",
        2912 => x"01010100",
        2913 => x"01010101",
        2914 => x"01010101",
        2915 => x"01010101",
        2916 => x"01010101",
        2917 => x"01000101",
        2918 => x"01000101",
        2919 => x"00010101",
        2920 => x"01010101",
        2921 => x"01010101",
        2922 => x"01010101",
        2923 => x"01010101",
        2924 => x"01010101",
        2925 => x"01010101",
        2926 => x"01010101",
        2927 => x"01010101",
        2928 => x"01010101",
        2929 => x"01010101",
        2930 => x"02010101",
        2931 => x"01010101",
        2932 => x"01010101",
        2933 => x"00010101",
        2934 => x"02020101",
        2935 => x"00010100",
        2936 => x"01010101",
        2937 => x"01010101",
        2938 => x"01010101",
        2939 => x"01010101",
        2940 => x"01010101",
        2941 => x"01010101",
        2942 => x"01010101",

                --  sprite 42
        2943 => x"03030300",
        2944 => x"03030303",
        2945 => x"01010101",
        2946 => x"01010101",
        2947 => x"03030303",
        2948 => x"03030101",
        2949 => x"01010101",
        2950 => x"01010101",
        2951 => x"03030303",
        2952 => x"03010101",
        2953 => x"01010101",
        2954 => x"01010101",
        2955 => x"03000301",
        2956 => x"01010101",
        2957 => x"01010101",
        2958 => x"01010101",
        2959 => x"03030302",
        2960 => x"01010101",
        2961 => x"01010101",
        2962 => x"01010101",
        2963 => x"03030302",
        2964 => x"02010101",
        2965 => x"01010101",
        2966 => x"01010101",
        2967 => x"03030302",
        2968 => x"01010101",
        2969 => x"01010101",
        2970 => x"01010101",
        2971 => x"00030301",
        2972 => x"01010101",
        2973 => x"01010101",
        2974 => x"01010101",
        2975 => x"03010101",
        2976 => x"01010101",
        2977 => x"01010101",
        2978 => x"01010101",
        2979 => x"03010101",
        2980 => x"01010101",
        2981 => x"01010101",
        2982 => x"01010101",
        2983 => x"03010101",
        2984 => x"01010101",
        2985 => x"01010101",
        2986 => x"01010101",
        2987 => x"01010101",
        2988 => x"01010101",
        2989 => x"01010101",
        2990 => x"01010101",
        2991 => x"01010101",
        2992 => x"01010101",
        2993 => x"01010101",
        2994 => x"01010101",
        2995 => x"01010101",
        2996 => x"01010101",
        2997 => x"01010101",
        2998 => x"01010101",
        2999 => x"01010101",
        3000 => x"01010101",
        3001 => x"01010101",
        3002 => x"01010101",
        3003 => x"01010101",
        3004 => x"01010101",
        3005 => x"01010101",
        3006 => x"01010101",

                --  sprite 43
        3007 => x"01010101",
        3008 => x"01010101",
        3009 => x"03030303",
        3010 => x"03000303",
        3011 => x"01010101",
        3012 => x"01010101",
        3013 => x"01030101",
        3014 => x"03030303",
        3015 => x"01010101",
        3016 => x"01010101",
        3017 => x"01010101",
        3018 => x"03030303",
        3019 => x"01010101",
        3020 => x"01010101",
        3021 => x"01010101",
        3022 => x"01010303",
        3023 => x"01010101",
        3024 => x"01010101",
        3025 => x"01010101",
        3026 => x"01010300",
        3027 => x"01010101",
        3028 => x"01010101",
        3029 => x"01010101",
        3030 => x"01010303",
        3031 => x"01010101",
        3032 => x"01010101",
        3033 => x"01010101",
        3034 => x"01010303",
        3035 => x"01010101",
        3036 => x"01010101",
        3037 => x"01010101",
        3038 => x"01010103",
        3039 => x"01010101",
        3040 => x"01010101",
        3041 => x"01010101",
        3042 => x"01010203",
        3043 => x"01010101",
        3044 => x"01010101",
        3045 => x"01010101",
        3046 => x"01020203",
        3047 => x"01010101",
        3048 => x"01010101",
        3049 => x"01010101",
        3050 => x"01010101",
        3051 => x"01010101",
        3052 => x"01010101",
        3053 => x"01010101",
        3054 => x"01010101",
        3055 => x"01010101",
        3056 => x"01010101",
        3057 => x"01010101",
        3058 => x"01010101",
        3059 => x"01010101",
        3060 => x"01010101",
        3061 => x"01010101",
        3062 => x"01010101",
        3063 => x"01010101",
        3064 => x"01010101",
        3065 => x"01010101",
        3066 => x"01010101",
        3067 => x"01010101",
        3068 => x"01010101",
        3069 => x"01010101",
        3070 => x"01010101",

                --  sprite 44
        3071 => x"01010101",
        3072 => x"01010101",
        3073 => x"01010101",
        3074 => x"01010101",
        3075 => x"01010101",
        3076 => x"01010101",
        3077 => x"01010101",
        3078 => x"01010101",
        3079 => x"01010101",
        3080 => x"01010101",
        3081 => x"01010101",
        3082 => x"01010101",
        3083 => x"01010101",
        3084 => x"01010101",
        3085 => x"01010101",
        3086 => x"01010101",
        3087 => x"02010101",
        3088 => x"01010101",
        3089 => x"01010101",
        3090 => x"01010101",
        3091 => x"02010101",
        3092 => x"01010101",
        3093 => x"01010101",
        3094 => x"01010101",
        3095 => x"02010101",
        3096 => x"01010101",
        3097 => x"01010101",
        3098 => x"01010101",
        3099 => x"03020101",
        3100 => x"01010101",
        3101 => x"01010101",
        3102 => x"01010101",
        3103 => x"03020101",
        3104 => x"01010101",
        3105 => x"01010101",
        3106 => x"01010101",
        3107 => x"03020101",
        3108 => x"01010101",
        3109 => x"01010101",
        3110 => x"01010101",
        3111 => x"03020101",
        3112 => x"01010101",
        3113 => x"01010101",
        3114 => x"01010101",
        3115 => x"00030202",
        3116 => x"01010101",
        3117 => x"01010101",
        3118 => x"01010101",
        3119 => x"03030302",
        3120 => x"01010101",
        3121 => x"01010101",
        3122 => x"01010101",
        3123 => x"03030302",
        3124 => x"02020101",
        3125 => x"01010101",
        3126 => x"01010101",
        3127 => x"03000302",
        3128 => x"02020201",
        3129 => x"01010101",
        3130 => x"01010101",
        3131 => x"03030303",
        3132 => x"03030202",
        3133 => x"01010101",
        3134 => x"01010101",

                --  sprite 45
        3135 => x"01010101",
        3136 => x"01010101",
        3137 => x"01010101",
        3138 => x"01010101",
        3139 => x"01010101",
        3140 => x"01010101",
        3141 => x"01010101",
        3142 => x"01010101",
        3143 => x"01010101",
        3144 => x"01010101",
        3145 => x"01010101",
        3146 => x"01010101",
        3147 => x"01010101",
        3148 => x"01010101",
        3149 => x"01010101",
        3150 => x"01010101",
        3151 => x"01010101",
        3152 => x"01010101",
        3153 => x"01010101",
        3154 => x"01010101",
        3155 => x"01010101",
        3156 => x"01010101",
        3157 => x"01010101",
        3158 => x"01010101",
        3159 => x"01010101",
        3160 => x"01010101",
        3161 => x"01010101",
        3162 => x"01010102",
        3163 => x"01010101",
        3164 => x"01010101",
        3165 => x"01010101",
        3166 => x"01010203",
        3167 => x"01010101",
        3168 => x"01010101",
        3169 => x"01010101",
        3170 => x"01010103",
        3171 => x"01010101",
        3172 => x"01010101",
        3173 => x"01010101",
        3174 => x"01010203",
        3175 => x"01010101",
        3176 => x"01010101",
        3177 => x"01010101",
        3178 => x"01020303",
        3179 => x"01010101",
        3180 => x"01010101",
        3181 => x"01010101",
        3182 => x"01020300",
        3183 => x"01010101",
        3184 => x"01010101",
        3185 => x"01010101",
        3186 => x"01020303",
        3187 => x"01010101",
        3188 => x"01010101",
        3189 => x"01010202",
        3190 => x"02030303",
        3191 => x"01010101",
        3192 => x"01010101",
        3193 => x"01010102",
        3194 => x"02030303",
        3195 => x"01010101",
        3196 => x"01010101",
        3197 => x"02020203",
        3198 => x"03030300",

                --  sprite 46
        3199 => x"03010303",
        3200 => x"03030303",
        3201 => x"00030302",
        3202 => x"03030303",
        3203 => x"03010303",
        3204 => x"03020303",
        3205 => x"00030302",
        3206 => x"03000303",
        3207 => x"01010303",
        3208 => x"01020303",
        3209 => x"00000303",
        3210 => x"03000301",
        3211 => x"00000303",
        3212 => x"01030103",
        3213 => x"00010300",
        3214 => x"03010101",
        3215 => x"01000103",
        3216 => x"00010103",
        3217 => x"01000301",
        3218 => x"03030100",
        3219 => x"01000101",
        3220 => x"01010001",
        3221 => x"01000101",
        3222 => x"03010100",
        3223 => x"01010103",
        3224 => x"01010101",
        3225 => x"01030101",
        3226 => x"03030301",
        3227 => x"01030103",
        3228 => x"01010301",
        3229 => x"03030103",
        3230 => x"03010301",
        3231 => x"03030103",
        3232 => x"03010301",
        3233 => x"03020302",
        3234 => x"03010301",
        3235 => x"03030303",
        3236 => x"03030301",
        3237 => x"03020303",
        3238 => x"03010303",
        3239 => x"03030302",
        3240 => x"03010303",
        3241 => x"03020303",
        3242 => x"03030303",
        3243 => x"03030302",
        3244 => x"03010303",
        3245 => x"03030303",
        3246 => x"03030303",
        3247 => x"03030103",
        3248 => x"03010303",
        3249 => x"03030303",
        3250 => x"03030303",
        3251 => x"03030303",
        3252 => x"03030303",
        3253 => x"01030303",
        3254 => x"03030301",
        3255 => x"03030303",
        3256 => x"03030303",
        3257 => x"03030303",
        3258 => x"03030303",
        3259 => x"03030303",
        3260 => x"03030303",
        3261 => x"03030303",
        3262 => x"03030303",

                --  sprite 47
        3263 => x"00000000",
        3264 => x"00000003",
        3265 => x"00000000",
        3266 => x"00000003",
        3267 => x"00020000",
        3268 => x"00020002",
        3269 => x"00020000",
        3270 => x"00020002",
        3271 => x"00000000",
        3272 => x"00000002",
        3273 => x"00000000",
        3274 => x"00000002",
        3275 => x"00000000",
        3276 => x"00000002",
        3277 => x"00000000",
        3278 => x"00000002",
        3279 => x"00000000",
        3280 => x"00000002",
        3281 => x"00000000",
        3282 => x"00000002",
        3283 => x"00000000",
        3284 => x"00000002",
        3285 => x"00000000",
        3286 => x"00000002",
        3287 => x"00000000",
        3288 => x"00000002",
        3289 => x"00000000",
        3290 => x"00000002",
        3291 => x"00000000",
        3292 => x"00000002",
        3293 => x"00000000",
        3294 => x"00000002",
        3295 => x"00000000",
        3296 => x"00000002",
        3297 => x"00000000",
        3298 => x"00000002",
        3299 => x"00000000",
        3300 => x"00000002",
        3301 => x"00000000",
        3302 => x"00000002",
        3303 => x"00000000",
        3304 => x"00000002",
        3305 => x"00000000",
        3306 => x"00000002",
        3307 => x"00000000",
        3308 => x"00000002",
        3309 => x"00000000",
        3310 => x"00000002",
        3311 => x"00000000",
        3312 => x"00000002",
        3313 => x"00000000",
        3314 => x"00000002",
        3315 => x"00020000",
        3316 => x"00020002",
        3317 => x"00020000",
        3318 => x"00020002",
        3319 => x"00000000",
        3320 => x"00000002",
        3321 => x"00000000",
        3322 => x"00000002",
        3323 => x"03020202",
        3324 => x"02020202",
        3325 => x"03020202",
        3326 => x"02020202",

                --  sprite 48
        3327 => x"01010101",
        3328 => x"01010101",
        3329 => x"01010101",
        3330 => x"01010101",
        3331 => x"01010101",
        3332 => x"01030303",
        3333 => x"03030301",
        3334 => x"01010103",
        3335 => x"02010103",
        3336 => x"03000000",
        3337 => x"00000002",
        3338 => x"02010103",
        3339 => x"02010300",
        3340 => x"00000000",
        3341 => x"00000000",
        3342 => x"00020103",
        3343 => x"02010300",
        3344 => x"00030303",
        3345 => x"03030300",
        3346 => x"00020103",
        3347 => x"00030000",
        3348 => x"03000202",
        3349 => x"02020002",
        3350 => x"00000200",
        3351 => x"00000003",
        3352 => x"00000202",
        3353 => x"02020000",
        3354 => x"02000000",
        3355 => x"00000003",
        3356 => x"00000000",
        3357 => x"00000000",
        3358 => x"02000000",
        3359 => x"00000003",
        3360 => x"00000303",
        3361 => x"03030000",
        3362 => x"02000000",
        3363 => x"00000000",
        3364 => x"02030200",
        3365 => x"00020302",
        3366 => x"00000000",
        3367 => x"00000000",
        3368 => x"03000200",
        3369 => x"00020003",
        3370 => x"00000000",
        3371 => x"00000101",
        3372 => x"01010100",
        3373 => x"00010101",
        3374 => x"01010000",
        3375 => x"00010000",
        3376 => x"02000001",
        3377 => x"01000002",
        3378 => x"00000100",
        3379 => x"01020000",
        3380 => x"02020002",
        3381 => x"02000202",
        3382 => x"00000201",
        3383 => x"01020200",
        3384 => x"02020202",
        3385 => x"02020202",
        3386 => x"00020201",
        3387 => x"02020200",
        3388 => x"02020202",
        3389 => x"02020202",
        3390 => x"00020202",

                --  sprite 49
        3391 => x"03010303",
        3392 => x"03030303",
        3393 => x"00030302",
        3394 => x"03030303",
        3395 => x"03010303",
        3396 => x"03020303",
        3397 => x"00030302",
        3398 => x"03000303",
        3399 => x"01010303",
        3400 => x"01020303",
        3401 => x"00000303",
        3402 => x"03000301",
        3403 => x"00000303",
        3404 => x"01030103",
        3405 => x"00010300",
        3406 => x"03010101",
        3407 => x"01000103",
        3408 => x"00010103",
        3409 => x"01000301",
        3410 => x"03030100",
        3411 => x"01000101",
        3412 => x"01010001",
        3413 => x"01000101",
        3414 => x"03010100",
        3415 => x"01010103",
        3416 => x"01010101",
        3417 => x"01030101",
        3418 => x"03030301",
        3419 => x"01030103",
        3420 => x"01010301",
        3421 => x"03030103",
        3422 => x"03010301",
        3423 => x"03030303",
        3424 => x"03030300",
        3425 => x"03030303",
        3426 => x"03030300",
        3427 => x"03030303",
        3428 => x"03030303",
        3429 => x"03030303",
        3430 => x"03030303",
        3431 => x"00030303",
        3432 => x"03030303",
        3433 => x"00030303",
        3434 => x"03030303",
        3435 => x"03030303",
        3436 => x"03030303",
        3437 => x"03030303",
        3438 => x"03030303",
        3439 => x"03030303",
        3440 => x"03030303",
        3441 => x"03030303",
        3442 => x"03030303",
        3443 => x"03030303",
        3444 => x"03030303",
        3445 => x"03030303",
        3446 => x"03030303",
        3447 => x"00030300",
        3448 => x"03010303",
        3449 => x"00030300",
        3450 => x"03010303",
        3451 => x"03030103",
        3452 => x"01010101",
        3453 => x"03030103",
        3454 => x"01010101",

                --  sprite 50
        3455 => x"06060606",
        3456 => x"06060505",
        3457 => x"05060606",
        3458 => x"06060606",
        3459 => x"06060606",
        3460 => x"06050505",
        3461 => x"05030606",
        3462 => x"06060606",
        3463 => x"06060606",
        3464 => x"05050505",
        3465 => x"05050306",
        3466 => x"06060606",
        3467 => x"06060605",
        3468 => x"05050303",
        3469 => x"02050503",
        3470 => x"06060606",
        3471 => x"06060505",
        3472 => x"05050303",
        3473 => x"02050505",
        3474 => x"03060606",
        3475 => x"06060505",
        3476 => x"03030303",
        3477 => x"03030205",
        3478 => x"03060606",
        3479 => x"06060505",
        3480 => x"03030303",
        3481 => x"03030205",
        3482 => x"03060606",
        3483 => x"06060505",
        3484 => x"02020303",
        3485 => x"02020205",
        3486 => x"03060606",
        3487 => x"03030505",
        3488 => x"05050303",
        3489 => x"02050505",
        3490 => x"03030306",
        3491 => x"03020505",
        3492 => x"05050303",
        3493 => x"02050505",
        3494 => x"03020302",
        3495 => x"03020505",
        3496 => x"05050502",
        3497 => x"02050505",
        3498 => x"03020302",
        3499 => x"03020505",
        3500 => x"05050505",
        3501 => x"05050505",
        3502 => x"03020302",
        3503 => x"03030303",
        3504 => x"03030303",
        3505 => x"03030303",
        3506 => x"03030302",
        3507 => x"05050505",
        3508 => x"05050505",
        3509 => x"05050505",
        3510 => x"05050502",
        3511 => x"05050505",
        3512 => x"05050505",
        3513 => x"05050505",
        3514 => x"05050502",
        3515 => x"02020202",
        3516 => x"02020202",
        3517 => x"02020202",
        3518 => x"02020202",

--			ENEMIES SPRITES
		        --  sprite 0
        4596 => x"00000000",		-- 35, 35, 35, 35
        4597 => x"00000000",		-- 35, 35, 35, 35
        4598 => x"00000000",		-- 35, 35, 35, 35
        4599 => x"00000000",		-- 35, 35, 35, 35
        4600 => x"00000000",		-- 35, 35, 35, 35
        4601 => x"00242428",		-- 35, 36, 36, 40
        4602 => x"28242400",		-- 40, 36, 36, 35
        4603 => x"00000000",		-- 35, 35, 35, 35
        4604 => x"24240024",		-- 36, 36, 35, 36
        4605 => x"24282424",		-- 36, 40, 36, 36
        4606 => x"24242824",		-- 36, 36, 40, 36
        4607 => x"24002424",		-- 36, 35, 36, 36
        4608 => x"00242424",		-- 35, 36, 36, 36
        4609 => x"24242424",		-- 36, 36, 36, 36
        4610 => x"24242424",		-- 36, 36, 36, 36
        4611 => x"24242400",		-- 36, 36, 36, 35
        4612 => x"00002424",		-- 35, 35, 36, 36
        4613 => x"24242824",		-- 36, 36, 40, 36
        4614 => x"24282424",		-- 36, 40, 36, 36
        4615 => x"24240000",		-- 36, 36, 35, 35
        4616 => x"24242424",		-- 36, 36, 36, 36
        4617 => x"28242424",		-- 40, 36, 36, 36
        4618 => x"24242428",		-- 36, 36, 36, 40
        4619 => x"24242424",		-- 36, 36, 36, 36
        4620 => x"00242424",		-- 35, 36, 36, 36
        4621 => x"27272424",		-- 39, 39, 36, 36
        4622 => x"24242727",		-- 36, 36, 39, 39
        4623 => x"24242400",		-- 36, 36, 36, 35
        4624 => x"00002427",		-- 35, 35, 36, 39
        4625 => x"27242727",		-- 39, 36, 39, 39
        4626 => x"27272427",		-- 39, 39, 36, 39
        4627 => x"27240000",		-- 39, 36, 35, 35
        4628 => x"00242427",		-- 35, 36, 36, 39
        4629 => x"27242427",		-- 39, 36, 36, 39
        4630 => x"27242427",		-- 39, 36, 36, 39
        4631 => x"27242400",		-- 39, 36, 36, 35
        4632 => x"24242424",		-- 36, 36, 36, 36
        4633 => x"27242427",		-- 39, 36, 36, 39
        4634 => x"27242427",		-- 39, 36, 36, 39
        4635 => x"24242424",		-- 36, 36, 36, 36
        4636 => x"00000024",		-- 35, 35, 35, 36
        4637 => x"27272427",		-- 39, 39, 36, 39
        4638 => x"27242727",		-- 39, 36, 39, 39
        4639 => x"24000000",		-- 36, 35, 35, 35
        4640 => x"00000024",		-- 35, 35, 35, 36
        4641 => x"24242727",		-- 36, 36, 39, 39
        4642 => x"27272424",		-- 39, 39, 36, 36
        4643 => x"24000000",		-- 36, 35, 35, 35
        4644 => x"00002424",		-- 35, 35, 36, 36
        4645 => x"00002424",		-- 35, 35, 36, 36
        4646 => x"24240000",		-- 36, 36, 35, 35
        4647 => x"24240000",		-- 36, 36, 35, 35
        4648 => x"00000000",		-- 35, 35, 35, 35
        4649 => x"00242424",		-- 35, 36, 36, 36
        4650 => x"24242400",		-- 36, 36, 36, 35
        4651 => x"00000000",		-- 35, 35, 35, 35
        4652 => x"00000000",		-- 35, 35, 35, 35
        4653 => x"24242424",		-- 36, 36, 36, 36
        4654 => x"24242424",		-- 36, 36, 36, 36
        4655 => x"00000000",		-- 35, 35, 35, 35
        4656 => x"00000000",		-- 35, 35, 35, 35
        4657 => x"00000000",		-- 35, 35, 35, 35
        4658 => x"00000000",		-- 35, 35, 35, 35
        4659 => x"00000000",		-- 35, 35, 35, 35

                --  sprite 1
        4660 => x"00002400",		-- 35, 35, 36, 35
        4661 => x"00002400",		-- 35, 35, 36, 35
        4662 => x"00000000",		-- 35, 35, 35, 35
        4663 => x"00000000",		-- 35, 35, 35, 35
        4664 => x"00002400",		-- 35, 35, 36, 35
        4665 => x"00000024",		-- 35, 35, 35, 36
        4666 => x"00002400",		-- 35, 35, 36, 35
        4667 => x"28000000",		-- 40, 35, 35, 35
        4668 => x"00000000",		-- 35, 35, 35, 35
        4669 => x"00240024",		-- 35, 36, 35, 36
        4670 => x"24000024",		-- 36, 35, 35, 36
        4671 => x"00240000",		-- 35, 36, 35, 35
        4672 => x"00002800",		-- 35, 35, 40, 35
        4673 => x"00242424",		-- 35, 36, 36, 36
        4674 => x"24240024",		-- 36, 36, 35, 36
        4675 => x"00240000",		-- 35, 36, 35, 35
        4676 => x"00000024",		-- 35, 35, 35, 36
        4677 => x"00242424",		-- 35, 36, 36, 36
        4678 => x"24242424",		-- 36, 36, 36, 36
        4679 => x"00000000",		-- 35, 35, 35, 35
        4680 => x"00240024",		-- 35, 36, 35, 36
        4681 => x"24002424",		-- 36, 35, 36, 36
        4682 => x"24282424",		-- 36, 40, 36, 36
        4683 => x"00242800",		-- 35, 36, 40, 35
        4684 => x"00242424",		-- 35, 36, 36, 36
        4685 => x"24282424",		-- 36, 40, 36, 36
        4686 => x"24242824",		-- 36, 36, 40, 36
        4687 => x"24242400",		-- 36, 36, 36, 35
        4688 => x"24002424",		-- 36, 35, 36, 36
        4689 => x"24242424",		-- 36, 36, 36, 36
        4690 => x"28242824",		-- 40, 36, 40, 36
        4691 => x"24242400",		-- 36, 36, 36, 35
        4692 => x"24002424",		-- 36, 35, 36, 36
        4693 => x"24242824",		-- 36, 36, 40, 36
        4694 => x"28242828",		-- 40, 36, 40, 40
        4695 => x"24242400",		-- 36, 36, 36, 35
        4696 => x"24242424",		-- 36, 36, 36, 36
        4697 => x"24282428",		-- 36, 40, 36, 40
        4698 => x"28282828",		-- 40, 40, 40, 40
        4699 => x"28240024",		-- 40, 36, 35, 36
        4700 => x"24242424",		-- 36, 36, 36, 36
        4701 => x"28282828",		-- 40, 40, 40, 40
        4702 => x"27282824",		-- 39, 40, 40, 36
        4703 => x"28242424",		-- 40, 36, 36, 36
        4704 => x"00242428",		-- 35, 36, 36, 40
        4705 => x"28282728",		-- 40, 40, 39, 40
        4706 => x"27282728",		-- 39, 40, 39, 40
        4707 => x"28242424",		-- 40, 36, 36, 36
        4708 => x"00242428",		-- 35, 36, 36, 40
        4709 => x"28272727",		-- 40, 39, 39, 39
        4710 => x"27272828",		-- 39, 39, 40, 40
        4711 => x"24242400",		-- 36, 36, 36, 35
        4712 => x"00002424",		-- 35, 35, 36, 36
        4713 => x"28282727",		-- 40, 40, 39, 39
        4714 => x"27272828",		-- 39, 39, 40, 40
        4715 => x"24242400",		-- 36, 36, 36, 35
        4716 => x"00002424",		-- 35, 35, 36, 36
        4717 => x"24282828",		-- 36, 40, 40, 40
        4718 => x"28282424",		-- 40, 40, 36, 36
        4719 => x"24240000",		-- 36, 36, 35, 35
        4720 => x"00000000",		-- 35, 35, 35, 35
        4721 => x"24242424",		-- 36, 36, 36, 36
        4722 => x"24242400",		-- 36, 36, 36, 35
        4723 => x"00000000",		-- 35, 35, 35, 35

                --  sprite 2
        4724 => x"00000000",		-- 35, 35, 35, 35
        4725 => x"00000000",		-- 35, 35, 35, 35
        4726 => x"00000000",		-- 35, 35, 35, 35
        4727 => x"00000000",		-- 35, 35, 35, 35
        4728 => x"00000000",		-- 35, 35, 35, 35
        4729 => x"00000000",		-- 35, 35, 35, 35
        4730 => x"00000000",		-- 35, 35, 35, 35
        4731 => x"00000000",		-- 35, 35, 35, 35
        4732 => x"00000000",		-- 35, 35, 35, 35
        4733 => x"00000000",		-- 35, 35, 35, 35
        4734 => x"00000000",		-- 35, 35, 35, 35
        4735 => x"00000000",		-- 35, 35, 35, 35
        4736 => x"00000000",		-- 35, 35, 35, 35
        4737 => x"00002424",		-- 35, 35, 36, 36
        4738 => x"24240000",		-- 36, 36, 35, 35
        4739 => x"00000000",		-- 35, 35, 35, 35
        4740 => x"00000000",		-- 35, 35, 35, 35
        4741 => x"00242424",		-- 35, 36, 36, 36
        4742 => x"24242400",		-- 36, 36, 36, 35
        4743 => x"00000000",		-- 35, 35, 35, 35
        4744 => x"00000000",		-- 35, 35, 35, 35
        4745 => x"00242428",		-- 35, 36, 36, 40
        4746 => x"28242400",		-- 40, 36, 36, 35
        4747 => x"00000000",		-- 35, 35, 35, 35
        4748 => x"00000000",		-- 35, 35, 35, 35
        4749 => x"24242828",		-- 36, 36, 40, 40
        4750 => x"28282424",		-- 40, 40, 36, 36
        4751 => x"00000000",		-- 35, 35, 35, 35
        4752 => x"00000000",		-- 35, 35, 35, 35
        4753 => x"24242827",		-- 36, 36, 40, 39
        4754 => x"27282424",		-- 39, 40, 36, 36
        4755 => x"00000000",		-- 35, 35, 35, 35
        4756 => x"00000000",		-- 35, 35, 35, 35
        4757 => x"24242827",		-- 36, 36, 40, 39
        4758 => x"27282424",		-- 39, 40, 36, 36
        4759 => x"00000000",		-- 35, 35, 35, 35
        4760 => x"00000000",		-- 35, 35, 35, 35
        4761 => x"24242828",		-- 36, 36, 40, 40
        4762 => x"28282424",		-- 40, 40, 36, 36
        4763 => x"00000000",		-- 35, 35, 35, 35
        4764 => x"00000000",		-- 35, 35, 35, 35
        4765 => x"00242428",		-- 35, 36, 36, 40
        4766 => x"28242400",		-- 40, 36, 36, 35
        4767 => x"00000000",		-- 35, 35, 35, 35
        4768 => x"00000000",		-- 35, 35, 35, 35
        4769 => x"00242424",		-- 35, 36, 36, 36
        4770 => x"24242400",		-- 36, 36, 36, 35
        4771 => x"00000000",		-- 35, 35, 35, 35
        4772 => x"00000000",		-- 35, 35, 35, 35
        4773 => x"00002424",		-- 35, 35, 36, 36
        4774 => x"24240000",		-- 36, 36, 35, 35
        4775 => x"00000000",		-- 35, 35, 35, 35
        4776 => x"00000000",		-- 35, 35, 35, 35
        4777 => x"00000000",		-- 35, 35, 35, 35
        4778 => x"00000000",		-- 35, 35, 35, 35
        4779 => x"00000000",		-- 35, 35, 35, 35
        4780 => x"00000000",		-- 35, 35, 35, 35
        4781 => x"00000000",		-- 35, 35, 35, 35
        4782 => x"00000000",		-- 35, 35, 35, 35
        4783 => x"00000000",		-- 35, 35, 35, 35
        4784 => x"00000000",		-- 35, 35, 35, 35
        4785 => x"00000000",		-- 35, 35, 35, 35
        4786 => x"00000000",		-- 35, 35, 35, 35
        4787 => x"00000000",		-- 35, 35, 35, 35

                --  sprite 3
        4788 => x"00000000",		-- 35, 35, 35, 35
        4789 => x"00242428",		-- 35, 36, 36, 40
        4790 => x"28242400",		-- 40, 36, 36, 35
        4791 => x"00000000",		-- 35, 35, 35, 35
        4792 => x"00000024",		-- 35, 35, 35, 36
        4793 => x"24282424",		-- 36, 40, 36, 36
        4794 => x"24242824",		-- 36, 36, 40, 36
        4795 => x"24000000",		-- 36, 35, 35, 35
        4796 => x"24242424",		-- 36, 36, 36, 36
        4797 => x"24242424",		-- 36, 36, 36, 36
        4798 => x"24242424",		-- 36, 36, 36, 36
        4799 => x"24242424",		-- 36, 36, 36, 36
        4800 => x"00242424",		-- 35, 36, 36, 36
        4801 => x"24242824",		-- 36, 36, 40, 36
        4802 => x"24282424",		-- 36, 40, 36, 36
        4803 => x"24242400",		-- 36, 36, 36, 35
        4804 => x"00002424",		-- 35, 35, 36, 36
        4805 => x"28242424",		-- 40, 36, 36, 36
        4806 => x"24242428",		-- 36, 36, 36, 40
        4807 => x"24240000",		-- 36, 36, 35, 35
        4808 => x"24242424",		-- 36, 36, 36, 36
        4809 => x"27272424",		-- 39, 39, 36, 36
        4810 => x"24242727",		-- 36, 36, 39, 39
        4811 => x"24242424",		-- 36, 36, 36, 36
        4812 => x"00242427",		-- 35, 36, 36, 39
        4813 => x"27242727",		-- 39, 36, 39, 39
        4814 => x"27272427",		-- 39, 39, 36, 39
        4815 => x"27242400",		-- 39, 36, 36, 35
        4816 => x"00002427",		-- 35, 35, 36, 39
        4817 => x"27242427",		-- 39, 36, 36, 39
        4818 => x"27242427",		-- 39, 36, 36, 39
        4819 => x"27240000",		-- 39, 36, 35, 35
        4820 => x"00242424",		-- 35, 36, 36, 36
        4821 => x"27242427",		-- 39, 36, 36, 39
        4822 => x"27242427",		-- 39, 36, 36, 39
        4823 => x"24242400",		-- 36, 36, 36, 35
        4824 => x"00240024",		-- 35, 36, 35, 36
        4825 => x"27272427",		-- 39, 39, 36, 39
        4826 => x"27242727",		-- 39, 36, 39, 39
        4827 => x"24002400",		-- 36, 35, 36, 35
        4828 => x"00000024",		-- 35, 35, 35, 36
        4829 => x"24242727",		-- 36, 36, 39, 39
        4830 => x"27272424",		-- 39, 39, 36, 36
        4831 => x"24000000",		-- 36, 35, 35, 35
        4832 => x"00000024",		-- 35, 35, 35, 36
        4833 => x"24002424",		-- 36, 35, 36, 36
        4834 => x"24240024",		-- 36, 36, 35, 36
        4835 => x"24000000",		-- 36, 35, 35, 35
        4836 => x"00000000",		-- 35, 35, 35, 35
        4837 => x"00002424",		-- 35, 35, 36, 36
        4838 => x"24240000",		-- 36, 36, 35, 35
        4839 => x"00000000",		-- 35, 35, 35, 35
        4840 => x"00000000",		-- 35, 35, 35, 35
        4841 => x"00002424",		-- 35, 35, 36, 36
        4842 => x"24240000",		-- 36, 36, 35, 35
        4843 => x"00000000",		-- 35, 35, 35, 35
        4844 => x"00000000",		-- 35, 35, 35, 35
        4845 => x"00002424",		-- 35, 35, 36, 36
        4846 => x"24240000",		-- 36, 36, 35, 35
        4847 => x"00000000",		-- 35, 35, 35, 35
        4848 => x"00000000",		-- 35, 35, 35, 35
        4849 => x"24242424",		-- 36, 36, 36, 36
        4850 => x"24242424",		-- 36, 36, 36, 36
        4851 => x"00000000",		-- 35, 35, 35, 35

                --  sprite 4
        4852 => x"00000000",		-- 35, 35, 35, 35
        4853 => x"00000000",		-- 35, 35, 35, 35
        4854 => x"00240000",		-- 35, 36, 35, 35
        4855 => x"00240000",		-- 35, 36, 35, 35
        4856 => x"00000028",		-- 35, 35, 35, 40
        4857 => x"00240000",		-- 35, 36, 35, 35
        4858 => x"24000000",		-- 36, 35, 35, 35
        4859 => x"00240000",		-- 35, 36, 35, 35
        4860 => x"00002400",		-- 35, 35, 36, 35
        4861 => x"24000024",		-- 36, 35, 35, 36
        4862 => x"24002400",		-- 36, 35, 36, 35
        4863 => x"00000000",		-- 35, 35, 35, 35
        4864 => x"00002400",		-- 35, 35, 36, 35
        4865 => x"24002424",		-- 36, 35, 36, 36
        4866 => x"24242400",		-- 36, 36, 36, 35
        4867 => x"00280000",		-- 35, 40, 35, 35
        4868 => x"00000000",		-- 35, 35, 35, 35
        4869 => x"24242424",		-- 36, 36, 36, 36
        4870 => x"24242400",		-- 36, 36, 36, 35
        4871 => x"24000000",		-- 36, 35, 35, 35
        4872 => x"00282400",		-- 35, 40, 36, 35
        4873 => x"24242824",		-- 36, 36, 40, 36
        4874 => x"24240024",		-- 36, 36, 35, 36
        4875 => x"24002400",		-- 36, 35, 36, 35
        4876 => x"00242424",		-- 35, 36, 36, 36
        4877 => x"24282424",		-- 36, 40, 36, 36
        4878 => x"24242824",		-- 36, 36, 40, 36
        4879 => x"24242400",		-- 36, 36, 36, 35
        4880 => x"00242424",		-- 35, 36, 36, 36
        4881 => x"24282428",		-- 36, 40, 36, 40
        4882 => x"24242424",		-- 36, 36, 36, 36
        4883 => x"24240024",		-- 36, 36, 35, 36
        4884 => x"00242424",		-- 35, 36, 36, 36
        4885 => x"28282428",		-- 40, 40, 36, 40
        4886 => x"24282424",		-- 36, 40, 36, 36
        4887 => x"24240024",		-- 36, 36, 35, 36
        4888 => x"24002428",		-- 36, 35, 36, 40
        4889 => x"28282828",		-- 40, 40, 40, 40
        4890 => x"28242824",		-- 40, 36, 40, 36
        4891 => x"24242424",		-- 36, 36, 36, 36
        4892 => x"24242428",		-- 36, 36, 36, 40
        4893 => x"24282827",		-- 36, 40, 40, 39
        4894 => x"28282828",		-- 40, 40, 40, 40
        4895 => x"24242424",		-- 36, 36, 36, 36
        4896 => x"24242428",		-- 36, 36, 36, 40
        4897 => x"28272827",		-- 40, 39, 40, 39
        4898 => x"28272828",		-- 40, 39, 40, 40
        4899 => x"28242400",		-- 40, 36, 36, 35
        4900 => x"00242424",		-- 35, 36, 36, 36
        4901 => x"28282727",		-- 40, 40, 39, 39
        4902 => x"27272728",		-- 39, 39, 39, 40
        4903 => x"28242400",		-- 40, 36, 36, 35
        4904 => x"00242424",		-- 35, 36, 36, 36
        4905 => x"28282727",		-- 40, 40, 39, 39
        4906 => x"27272828",		-- 39, 39, 40, 40
        4907 => x"24240000",		-- 36, 36, 35, 35
        4908 => x"00002424",		-- 35, 35, 36, 36
        4909 => x"24242828",		-- 36, 36, 40, 40
        4910 => x"28282824",		-- 40, 40, 40, 36
        4911 => x"24240000",		-- 36, 36, 35, 35
        4912 => x"00000000",		-- 35, 35, 35, 35
        4913 => x"00242424",		-- 35, 36, 36, 36
        4914 => x"24242424",		-- 36, 36, 36, 36
        4915 => x"00000000",		-- 35, 35, 35, 35

                --  sprite 5
        4916 => x"00000000",		-- 35, 35, 35, 35
        4917 => x"00272727",		-- 35, 39, 39, 39
        4918 => x"27272700",		-- 39, 39, 39, 35
        4919 => x"00000000",		-- 35, 35, 35, 35
        4920 => x"27000026",		-- 39, 35, 35, 38
        4921 => x"26262626",		-- 38, 38, 38, 38
        4922 => x"25272727",		-- 37, 39, 39, 39
        4923 => x"26000000",		-- 38, 35, 35, 35
        4924 => x"27002626",		-- 39, 35, 38, 38
        4925 => x"25252626",		-- 37, 37, 38, 38
        4926 => x"26252726",		-- 38, 37, 39, 38
        4927 => x"00002726",		-- 35, 35, 39, 38
        4928 => x"27272625",		-- 39, 39, 38, 37
        4929 => x"25252526",		-- 37, 37, 37, 38
        4930 => x"25272626",		-- 37, 39, 38, 38
        4931 => x"27272600",		-- 39, 39, 38, 35
        4932 => x"27272727",		-- 39, 39, 39, 39
        4933 => x"27272727",		-- 39, 39, 39, 39
        4934 => x"27272727",		-- 39, 39, 39, 39
        4935 => x"27260000",		-- 39, 38, 35, 35
        4936 => x"00272526",		-- 35, 39, 37, 38
        4937 => x"26262525",		-- 38, 38, 37, 37
        4938 => x"27272727",		-- 39, 39, 39, 39
        4939 => x"26000000",		-- 38, 35, 35, 35
        4940 => x"00252525",		-- 35, 37, 37, 37
        4941 => x"25252525",		-- 37, 37, 37, 37
        4942 => x"25272726",		-- 37, 39, 39, 38
        4943 => x"26000000",		-- 38, 35, 35, 35
        4944 => x"00252525",		-- 35, 37, 37, 37
        4945 => x"25252525",		-- 37, 37, 37, 37
        4946 => x"25252726",		-- 37, 37, 39, 38
        4947 => x"00000000",		-- 35, 35, 35, 35
        4948 => x"00252527",		-- 35, 37, 37, 39
        4949 => x"27272525",		-- 39, 39, 37, 37
        4950 => x"25252726",		-- 37, 37, 39, 38
        4951 => x"00000000",		-- 35, 35, 35, 35
        4952 => x"00002727",		-- 35, 35, 39, 39
        4953 => x"27272727",		-- 39, 39, 39, 39
        4954 => x"27272726",		-- 39, 39, 39, 38
        4955 => x"00000000",		-- 35, 35, 35, 35
        4956 => x"00000027",		-- 35, 35, 35, 39
        4957 => x"27272727",		-- 39, 39, 39, 39
        4958 => x"27272727",		-- 39, 39, 39, 39
        4959 => x"26000000",		-- 38, 35, 35, 35
        4960 => x"00000000",		-- 35, 35, 35, 35
        4961 => x"27272727",		-- 39, 39, 39, 39
        4962 => x"27272727",		-- 39, 39, 39, 39
        4963 => x"26000000",		-- 38, 35, 35, 35
        4964 => x"00000000",		-- 35, 35, 35, 35
        4965 => x"00002727",		-- 35, 35, 39, 39
        4966 => x"27272727",		-- 39, 39, 39, 39
        4967 => x"27260000",		-- 39, 38, 35, 35
        4968 => x"00000025",		-- 35, 35, 35, 37
        4969 => x"25252525",		-- 37, 37, 37, 37
        4970 => x"25252727",		-- 37, 37, 39, 39
        4971 => x"27272600",		-- 39, 39, 38, 35
        4972 => x"00002525",		-- 35, 35, 37, 37
        4973 => x"25252525",		-- 37, 37, 37, 37
        4974 => x"25252525",		-- 37, 37, 37, 37
        4975 => x"25252525",		-- 37, 37, 37, 37
        4976 => x"00000000",		-- 35, 35, 35, 35
        4977 => x"25252525",		-- 37, 37, 37, 37
        4978 => x"25252525",		-- 37, 37, 37, 37
        4979 => x"25252500",		-- 37, 37, 37, 35

                --  sprite 6
        4980 => x"00000000",		-- 35, 35, 35, 35
        4981 => x"00272727",		-- 35, 39, 39, 39
        4982 => x"27272700",		-- 39, 39, 39, 35
        4983 => x"00000000",		-- 35, 35, 35, 35
        4984 => x"00000026",		-- 35, 35, 35, 38
        4985 => x"27272725",		-- 39, 39, 39, 37
        4986 => x"26262626",		-- 38, 38, 38, 38
        4987 => x"26000027",		-- 38, 35, 35, 39
        4988 => x"26270000",		-- 38, 39, 35, 35
        4989 => x"26272526",		-- 38, 39, 37, 38
        4990 => x"26262525",		-- 38, 38, 37, 37
        4991 => x"26260027",		-- 38, 38, 35, 39
        4992 => x"00262727",		-- 35, 38, 39, 39
        4993 => x"26262725",		-- 38, 38, 39, 37
        4994 => x"26252525",		-- 38, 37, 37, 37
        4995 => x"25262727",		-- 37, 38, 39, 39
        4996 => x"00002627",		-- 35, 35, 38, 39
        4997 => x"27272727",		-- 39, 39, 39, 39
        4998 => x"27272727",		-- 39, 39, 39, 39
        4999 => x"27272727",		-- 39, 39, 39, 39
        5000 => x"00000026",		-- 35, 35, 35, 38
        5001 => x"27272727",		-- 39, 39, 39, 39
        5002 => x"25252626",		-- 37, 37, 38, 38
        5003 => x"26252700",		-- 38, 37, 39, 35
        5004 => x"00000026",		-- 35, 35, 35, 38
        5005 => x"26272725",		-- 38, 39, 39, 37
        5006 => x"25252525",		-- 37, 37, 37, 37
        5007 => x"25252500",		-- 37, 37, 37, 35
        5008 => x"00000000",		-- 35, 35, 35, 35
        5009 => x"26272525",		-- 38, 39, 37, 37
        5010 => x"25252525",		-- 37, 37, 37, 37
        5011 => x"25252500",		-- 37, 37, 37, 35
        5012 => x"00000000",		-- 35, 35, 35, 35
        5013 => x"26272525",		-- 38, 39, 37, 37
        5014 => x"25252727",		-- 37, 37, 39, 39
        5015 => x"27252500",		-- 39, 37, 37, 35
        5016 => x"00000000",		-- 35, 35, 35, 35
        5017 => x"26272727",		-- 38, 39, 39, 39
        5018 => x"27272727",		-- 39, 39, 39, 39
        5019 => x"27270000",		-- 39, 39, 35, 35
        5020 => x"00000026",		-- 35, 35, 35, 38
        5021 => x"27272727",		-- 39, 39, 39, 39
        5022 => x"27272727",		-- 39, 39, 39, 39
        5023 => x"27000000",		-- 39, 35, 35, 35
        5024 => x"00000026",		-- 35, 35, 35, 38
        5025 => x"27272727",		-- 39, 39, 39, 39
        5026 => x"27272727",		-- 39, 39, 39, 39
        5027 => x"00000000",		-- 35, 35, 35, 35
        5028 => x"00002627",		-- 35, 35, 38, 39
        5029 => x"27272727",		-- 39, 39, 39, 39
        5030 => x"27270000",		-- 39, 39, 35, 35
        5031 => x"00000000",		-- 35, 35, 35, 35
        5032 => x"00262727",		-- 35, 38, 39, 39
        5033 => x"27272525",		-- 39, 39, 37, 37
        5034 => x"25252525",		-- 37, 37, 37, 37
        5035 => x"25000000",		-- 37, 35, 35, 35
        5036 => x"25252525",		-- 37, 37, 37, 37
        5037 => x"25252525",		-- 37, 37, 37, 37
        5038 => x"25252525",		-- 37, 37, 37, 37
        5039 => x"25250000",		-- 37, 37, 35, 35
        5040 => x"00252525",		-- 35, 37, 37, 37
        5041 => x"25252525",		-- 37, 37, 37, 37
        5042 => x"25252525",		-- 37, 37, 37, 37
        5043 => x"00000000",		-- 35, 35, 35, 35

                --  sprite 7
        5044 => x"00000000",		-- 35, 35, 35, 35
        5045 => x"26262627",		-- 38, 38, 38, 39
        5046 => x"27270000",		-- 39, 39, 35, 35
        5047 => x"00000000",		-- 35, 35, 35, 35
        5048 => x"00000026",		-- 35, 35, 35, 38
        5049 => x"27272727",		-- 39, 39, 39, 39
        5050 => x"27272727",		-- 39, 39, 39, 39
        5051 => x"00000000",		-- 35, 35, 35, 35
        5052 => x"27272627",		-- 39, 39, 38, 39
        5053 => x"27272727",		-- 39, 39, 39, 39
        5054 => x"27272727",		-- 39, 39, 39, 39
        5055 => x"27002727",		-- 39, 35, 39, 39
        5056 => x"26272726",		-- 38, 39, 39, 38
        5057 => x"27272727",		-- 39, 39, 39, 39
        5058 => x"27272727",		-- 39, 39, 39, 39
        5059 => x"26272700",		-- 38, 39, 39, 35
        5060 => x"00262727",		-- 35, 38, 39, 39
        5061 => x"26272727",		-- 38, 39, 39, 39
        5062 => x"27272727",		-- 39, 39, 39, 39
        5063 => x"26272700",		-- 38, 39, 39, 35
        5064 => x"00002627",		-- 35, 35, 38, 39
        5065 => x"27272727",		-- 39, 39, 39, 39
        5066 => x"27272727",		-- 39, 39, 39, 39
        5067 => x"27270000",		-- 39, 39, 35, 35
        5068 => x"00002627",		-- 35, 35, 38, 39
        5069 => x"27272727",		-- 39, 39, 39, 39
        5070 => x"27272727",		-- 39, 39, 39, 39
        5071 => x"27260000",		-- 39, 38, 35, 35
        5072 => x"00000026",		-- 35, 35, 35, 38
        5073 => x"27272727",		-- 39, 39, 39, 39
        5074 => x"27272727",		-- 39, 39, 39, 39
        5075 => x"27000000",		-- 39, 35, 35, 35
        5076 => x"00000026",		-- 35, 35, 35, 38
        5077 => x"27272727",		-- 39, 39, 39, 39
        5078 => x"27272727",		-- 39, 39, 39, 39
        5079 => x"27000000",		-- 39, 35, 35, 35
        5080 => x"00000000",		-- 35, 35, 35, 35
        5081 => x"26272727",		-- 38, 39, 39, 39
        5082 => x"27272727",		-- 39, 39, 39, 39
        5083 => x"27270000",		-- 39, 39, 35, 35
        5084 => x"00000000",		-- 35, 35, 35, 35
        5085 => x"26272727",		-- 38, 39, 39, 39
        5086 => x"27272727",		-- 39, 39, 39, 39
        5087 => x"27270000",		-- 39, 39, 35, 35
        5088 => x"00000000",		-- 35, 35, 35, 35
        5089 => x"00262727",		-- 35, 38, 39, 39
        5090 => x"27272727",		-- 39, 39, 39, 39
        5091 => x"27272700",		-- 39, 39, 39, 35
        5092 => x"00000000",		-- 35, 35, 35, 35
        5093 => x"00002626",		-- 35, 35, 38, 38
        5094 => x"26272727",		-- 38, 39, 39, 39
        5095 => x"27272700",		-- 39, 39, 39, 35
        5096 => x"00000000",		-- 35, 35, 35, 35
        5097 => x"25252525",		-- 37, 37, 37, 37
        5098 => x"25262626",		-- 37, 38, 38, 38
        5099 => x"26272727",		-- 38, 39, 39, 39
        5100 => x"00000025",		-- 35, 35, 35, 37
        5101 => x"25252525",		-- 37, 37, 37, 37
        5102 => x"25252525",		-- 37, 37, 37, 37
        5103 => x"25252525",		-- 37, 37, 37, 37
        5104 => x"00000000",		-- 35, 35, 35, 35
        5105 => x"25252525",		-- 37, 37, 37, 37
        5106 => x"25252525",		-- 37, 37, 37, 37
        5107 => x"25252500",		-- 37, 37, 37, 35

                --  sprite 8
        5108 => x"00000000",		-- 35, 35, 35, 35
        5109 => x"00002727",		-- 35, 35, 39, 39
        5110 => x"27262626",		-- 39, 38, 38, 38
        5111 => x"00000000",		-- 35, 35, 35, 35
        5112 => x"00000000",		-- 35, 35, 35, 35
        5113 => x"27272727",		-- 39, 39, 39, 39
        5114 => x"27272727",		-- 39, 39, 39, 39
        5115 => x"26000000",		-- 38, 35, 35, 35
        5116 => x"27270027",		-- 39, 39, 35, 39
        5117 => x"27272727",		-- 39, 39, 39, 39
        5118 => x"27272727",		-- 39, 39, 39, 39
        5119 => x"27262727",		-- 39, 38, 39, 39
        5120 => x"00272726",		-- 35, 39, 39, 38
        5121 => x"27272727",		-- 39, 39, 39, 39
        5122 => x"27272727",		-- 39, 39, 39, 39
        5123 => x"26272726",		-- 38, 39, 39, 38
        5124 => x"00272726",		-- 35, 39, 39, 38
        5125 => x"27272727",		-- 39, 39, 39, 39
        5126 => x"27272726",		-- 39, 39, 39, 38
        5127 => x"27272600",		-- 39, 39, 38, 35
        5128 => x"00002727",		-- 35, 35, 39, 39
        5129 => x"27272727",		-- 39, 39, 39, 39
        5130 => x"27272727",		-- 39, 39, 39, 39
        5131 => x"27260000",		-- 39, 38, 35, 35
        5132 => x"00002627",		-- 35, 35, 38, 39
        5133 => x"27272727",		-- 39, 39, 39, 39
        5134 => x"27272727",		-- 39, 39, 39, 39
        5135 => x"27260000",		-- 39, 38, 35, 35
        5136 => x"00000027",		-- 35, 35, 35, 39
        5137 => x"27272727",		-- 39, 39, 39, 39
        5138 => x"27272727",		-- 39, 39, 39, 39
        5139 => x"26000000",		-- 38, 35, 35, 35
        5140 => x"00000027",		-- 35, 35, 35, 39
        5141 => x"27272727",		-- 39, 39, 39, 39
        5142 => x"27272727",		-- 39, 39, 39, 39
        5143 => x"26000000",		-- 38, 35, 35, 35
        5144 => x"00002727",		-- 35, 35, 39, 39
        5145 => x"27272727",		-- 39, 39, 39, 39
        5146 => x"27272726",		-- 39, 39, 39, 38
        5147 => x"00000000",		-- 35, 35, 35, 35
        5148 => x"00002727",		-- 35, 35, 39, 39
        5149 => x"27272727",		-- 39, 39, 39, 39
        5150 => x"27272726",		-- 39, 39, 39, 38
        5151 => x"00000000",		-- 35, 35, 35, 35
        5152 => x"00272727",		-- 35, 39, 39, 39
        5153 => x"27272727",		-- 39, 39, 39, 39
        5154 => x"27272600",		-- 39, 39, 38, 35
        5155 => x"00000000",		-- 35, 35, 35, 35
        5156 => x"00272727",		-- 35, 39, 39, 39
        5157 => x"27272726",		-- 39, 39, 39, 38
        5158 => x"26260000",		-- 38, 38, 35, 35
        5159 => x"00000000",		-- 35, 35, 35, 35
        5160 => x"27272726",		-- 39, 39, 39, 38
        5161 => x"26262625",		-- 38, 38, 38, 37
        5162 => x"25252525",		-- 37, 37, 37, 37
        5163 => x"00000000",		-- 35, 35, 35, 35
        5164 => x"25252525",		-- 37, 37, 37, 37
        5165 => x"25252525",		-- 37, 37, 37, 37
        5166 => x"25252525",		-- 37, 37, 37, 37
        5167 => x"25000000",		-- 37, 35, 35, 35
        5168 => x"00252525",		-- 35, 37, 37, 37
        5169 => x"25252525",		-- 37, 37, 37, 37
        5170 => x"25252525",		-- 37, 37, 37, 37
        5171 => x"00000000",		-- 35, 35, 35, 35
		
--          LINK SPRITES
                --  sprite 0
        5172 => x"00000000",		-- 8, 8, 8, 8
        5173 => x"00090909",		-- 8, 9, 9, 9
        5174 => x"09090900",		-- 9, 9, 9, 8
        5175 => x"00000000",		-- 8, 8, 8, 8
        5176 => x"00000000",		-- 8, 8, 8, 8
        5177 => x"09090909",		-- 9, 9, 9, 9
        5178 => x"09090909",		-- 9, 9, 9, 9
        5179 => x"00000000",		-- 8, 8, 8, 8
        5180 => x"00000A00",		-- 8, 8, 10, 8
        5181 => x"090B0B0B",		-- 9, 11, 11, 11
        5182 => x"0B0B0B09",		-- 11, 11, 11, 9
        5183 => x"000A0000",		-- 8, 10, 8, 8
        5184 => x"00000A00",		-- 8, 8, 10, 8
        5185 => x"0B0B0B0B",		-- 11, 11, 11, 11
        5186 => x"0B0B0B0B",		-- 11, 11, 11, 11
        5187 => x"000A0000",		-- 8, 10, 8, 8
        5188 => x"00000A0A",		-- 8, 8, 10, 10
        5189 => x"0B0A090A",		-- 11, 10, 9, 10
        5190 => x"0A090A0B",		-- 10, 9, 10, 11
        5191 => x"0A0A0000",		-- 10, 10, 8, 8
        5192 => x"00000A0A",		-- 8, 8, 10, 10
        5193 => x"0B0A0B0A",		-- 11, 10, 11, 10
        5194 => x"0A0B0A0B",		-- 10, 11, 10, 11
        5195 => x"0A0A0000",		-- 10, 10, 8, 8
        5196 => x"0000000A",		-- 8, 8, 8, 10
        5197 => x"0A0A0A0A",		-- 10, 10, 10, 10
        5198 => x"0A0A0A0A",		-- 10, 10, 10, 10
        5199 => x"0A0B0000",		-- 10, 11, 8, 8
        5200 => x"00000009",		-- 8, 8, 8, 9
        5201 => x"090A0A0B",		-- 9, 10, 10, 11
        5202 => x"0B0A0A09",		-- 11, 10, 10, 9
        5203 => x"090B0000",		-- 9, 11, 8, 8
        5204 => x"000B0B0B",		-- 8, 11, 11, 11
        5205 => x"0B0B0A0A",		-- 11, 11, 10, 10
        5206 => x"0A0A0909",		-- 10, 10, 9, 9
        5207 => x"0B0B0B00",		-- 11, 11, 11, 8
        5208 => x"0B0B0A0B",		-- 11, 11, 10, 11
        5209 => x"0B0B0B09",		-- 11, 11, 11, 9
        5210 => x"09090909",		-- 9, 9, 9, 9
        5211 => x"0A0B0B00",		-- 10, 11, 11, 8
        5212 => x"0B0A0A0A",		-- 11, 10, 10, 10
        5213 => x"0B0B0A0B",		-- 11, 11, 10, 11
        5214 => x"0B09090A",		-- 11, 9, 9, 10
        5215 => x"0A0A0B00",		-- 10, 10, 11, 8
        5216 => x"0B0B0A0B",		-- 11, 11, 10, 11
        5217 => x"0B0B0A09",		-- 11, 11, 10, 9
        5218 => x"0B0B0B0B",		-- 11, 11, 11, 11
        5219 => x"0A0A0A00",		-- 10, 10, 10, 8
        5220 => x"0B0B0A0B",		-- 11, 11, 10, 11
        5221 => x"0B0B0A0B",		-- 11, 11, 10, 11
        5222 => x"0B090909",		-- 11, 9, 9, 9
        5223 => x"090A0000",		-- 9, 10, 8, 8
        5224 => x"0B0B0B0B",		-- 11, 11, 11, 11
        5225 => x"0B0B0A09",		-- 11, 11, 10, 9
        5226 => x"09090909",		-- 9, 9, 9, 9
        5227 => x"00000000",		-- 8, 8, 8, 8
        5228 => x"000A0A0A",		-- 8, 10, 10, 10
        5229 => x"0A0A0B00",		-- 10, 10, 11, 8
        5230 => x"000B0B0B",		-- 8, 11, 11, 11
        5231 => x"00000000",		-- 8, 8, 8, 8
        5232 => x"00000000",		-- 8, 8, 8, 8
        5233 => x"0B0B0B00",		-- 11, 11, 11, 8
        5234 => x"00000000",		-- 8, 8, 8, 8
        5235 => x"00000000",		-- 8, 8, 8, 8

                --  sprite 1
        5236 => x"00000000",		-- 8, 8, 8, 8
        5237 => x"00090909",		-- 8, 9, 9, 9
        5238 => x"09090900",		-- 9, 9, 9, 8
        5239 => x"00000000",		-- 8, 8, 8, 8
        5240 => x"00000000",		-- 8, 8, 8, 8
        5241 => x"09090909",		-- 9, 9, 9, 9
        5242 => x"09090909",		-- 9, 9, 9, 9
        5243 => x"00000000",		-- 8, 8, 8, 8
        5244 => x"00000A00",		-- 8, 8, 10, 8
        5245 => x"090B0B0B",		-- 9, 11, 11, 11
        5246 => x"0B0B0B09",		-- 11, 11, 11, 9
        5247 => x"000A0000",		-- 8, 10, 8, 8
        5248 => x"00000A00",		-- 8, 8, 10, 8
        5249 => x"0B0B0B0B",		-- 11, 11, 11, 11
        5250 => x"0B0B0B0B",		-- 11, 11, 11, 11
        5251 => x"000A0000",		-- 8, 10, 8, 8
        5252 => x"00000A0A",		-- 8, 8, 10, 10
        5253 => x"0B0A090A",		-- 11, 10, 9, 10
        5254 => x"0A090A0B",		-- 10, 9, 10, 11
        5255 => x"0A0A0000",		-- 10, 10, 8, 8
        5256 => x"00000A0A",		-- 8, 8, 10, 10
        5257 => x"0B0A0B0A",		-- 11, 10, 11, 10
        5258 => x"0A0B0A0B",		-- 10, 11, 10, 11
        5259 => x"0A0A0000",		-- 10, 10, 8, 8
        5260 => x"0000000A",		-- 8, 8, 8, 10
        5261 => x"0A0A0A0A",		-- 10, 10, 10, 10
        5262 => x"0A0A0A0A",		-- 10, 10, 10, 10
        5263 => x"0A0B0000",		-- 10, 11, 8, 8
        5264 => x"00000000",		-- 8, 8, 8, 8
        5265 => x"090A0A0B",		-- 9, 10, 10, 11
        5266 => x"0B0A0A09",		-- 11, 10, 10, 9
        5267 => x"0B0B0000",		-- 11, 11, 8, 8
        5268 => x"00000B0B",		-- 8, 8, 11, 11
        5269 => x"0B0B0B0A",		-- 11, 11, 11, 10
        5270 => x"0A0A0909",		-- 10, 10, 9, 9
        5271 => x"090A0000",		-- 9, 10, 8, 8
        5272 => x"000B0B0A",		-- 8, 11, 11, 10
        5273 => x"0B0B0B0B",		-- 11, 11, 11, 11
        5274 => x"09090909",		-- 9, 9, 9, 9
        5275 => x"090A0000",		-- 9, 10, 8, 8
        5276 => x"000B0A0A",		-- 8, 11, 10, 10
        5277 => x"0A0B0B0A",		-- 10, 11, 11, 10
        5278 => x"0B0B0909",		-- 11, 11, 9, 9
        5279 => x"0B000000",		-- 11, 8, 8, 8
        5280 => x"000B0B0A",		-- 8, 11, 11, 10
        5281 => x"0B0B0B0A",		-- 11, 11, 11, 10
        5282 => x"090B0B0B",		-- 9, 11, 11, 11
        5283 => x"09000000",		-- 9, 8, 8, 8
        5284 => x"000B0B0A",		-- 8, 11, 11, 10
        5285 => x"0B0B0B0A",		-- 11, 11, 11, 10
        5286 => x"0B0B0909",		-- 11, 11, 9, 9
        5287 => x"09000000",		-- 9, 8, 8, 8
        5288 => x"000B0B0B",		-- 8, 11, 11, 11
        5289 => x"0B0B0B0A",		-- 11, 11, 11, 10
        5290 => x"0909090B",		-- 9, 9, 9, 11
        5291 => x"00000000",		-- 8, 8, 8, 8
        5292 => x"00000A0A",		-- 8, 8, 10, 10
        5293 => x"0A0A0A00",		-- 10, 10, 10, 8
        5294 => x"000B0B0B",		-- 8, 11, 11, 11
        5295 => x"00000000",		-- 8, 8, 8, 8
        5296 => x"00000000",		-- 8, 8, 8, 8
        5297 => x"00000000",		-- 8, 8, 8, 8
        5298 => x"000B0B0B",		-- 8, 11, 11, 11
        5299 => x"00000000",		-- 8, 8, 8, 8

                --  sprite 2
        5300 => x"00000000",		-- 8, 8, 8, 8
        5301 => x"00090909",		-- 8, 9, 9, 9
        5302 => x"09090900",		-- 9, 9, 9, 8
        5303 => x"00000000",		-- 8, 8, 8, 8
        5304 => x"00000000",		-- 8, 8, 8, 8
        5305 => x"09090909",		-- 9, 9, 9, 9
        5306 => x"09090909",		-- 9, 9, 9, 9
        5307 => x"00000000",		-- 8, 8, 8, 8
        5308 => x"00000A00",		-- 8, 8, 10, 8
        5309 => x"09090909",		-- 9, 9, 9, 9
        5310 => x"09090909",		-- 9, 9, 9, 9
        5311 => x"000A0000",		-- 8, 10, 8, 8
        5312 => x"00000A09",		-- 8, 8, 10, 9
        5313 => x"09090909",		-- 9, 9, 9, 9
        5314 => x"09090909",		-- 9, 9, 9, 9
        5315 => x"090A0000",		-- 9, 10, 8, 8
        5316 => x"00000A0B",		-- 8, 8, 10, 11
        5317 => x"09090909",		-- 9, 9, 9, 9
        5318 => x"09090909",		-- 9, 9, 9, 9
        5319 => x"0B0A0000",		-- 11, 10, 8, 8
        5320 => x"00000A0A",		-- 8, 8, 10, 10
        5321 => x"0B0B0909",		-- 11, 11, 9, 9
        5322 => x"09090B0B",		-- 9, 9, 11, 11
        5323 => x"0A0A0000",		-- 10, 10, 8, 8
        5324 => x"0000000A",		-- 8, 8, 8, 10
        5325 => x"0B0B0B09",		-- 11, 11, 11, 9
        5326 => x"090B0B0B",		-- 9, 11, 11, 11
        5327 => x"0A000000",		-- 10, 8, 8, 8
        5328 => x"0000000B",		-- 8, 8, 8, 11
        5329 => x"090B0B0B",		-- 9, 11, 11, 11
        5330 => x"0B0B0B09",		-- 11, 11, 11, 9
        5331 => x"0B000000",		-- 11, 8, 8, 8
        5332 => x"0000000B",		-- 8, 8, 8, 11
        5333 => x"0B090909",		-- 11, 9, 9, 9
        5334 => x"09090909",		-- 9, 9, 9, 9
        5335 => x"0B0B0000",		-- 11, 11, 8, 8
        5336 => x"00000A0B",		-- 8, 8, 10, 11
        5337 => x"0B090909",		-- 11, 9, 9, 9
        5338 => x"09090909",		-- 9, 9, 9, 9
        5339 => x"0B0B0000",		-- 11, 11, 8, 8
        5340 => x"00000A0B",		-- 8, 8, 10, 11
        5341 => x"0B090909",		-- 11, 9, 9, 9
        5342 => x"0909090B",		-- 9, 9, 9, 11
        5343 => x"0B000000",		-- 11, 8, 8, 8
        5344 => x"00000A0A",		-- 8, 8, 10, 10
        5345 => x"090B0B0B",		-- 9, 11, 11, 11
        5346 => x"0B0B0B09",		-- 11, 11, 11, 9
        5347 => x"09000000",		-- 9, 8, 8, 8
        5348 => x"00000009",		-- 8, 8, 8, 9
        5349 => x"09090909",		-- 9, 9, 9, 9
        5350 => x"09090909",		-- 9, 9, 9, 9
        5351 => x"09000000",		-- 9, 8, 8, 8
        5352 => x"00000000",		-- 8, 8, 8, 8
        5353 => x"0B090909",		-- 11, 9, 9, 9
        5354 => x"09090B0B",		-- 9, 9, 11, 11
        5355 => x"0B000000",		-- 11, 8, 8, 8
        5356 => x"00000000",		-- 8, 8, 8, 8
        5357 => x"000B0B00",		-- 8, 11, 11, 8
        5358 => x"000B0B0B",		-- 8, 11, 11, 11
        5359 => x"0B000000",		-- 11, 8, 8, 8
        5360 => x"00000000",		-- 8, 8, 8, 8
        5361 => x"00000000",		-- 8, 8, 8, 8
        5362 => x"00000B0B",		-- 8, 8, 11, 11
        5363 => x"00000000",		-- 8, 8, 8, 8

                --  sprite 3
        5364 => x"00000000",		-- 8, 8, 8, 8
        5365 => x"00000000",		-- 8, 8, 8, 8
        5366 => x"00000000",		-- 8, 8, 8, 8
        5367 => x"00000000",		-- 8, 8, 8, 8
        5368 => x"00000000",		-- 8, 8, 8, 8
        5369 => x"00090909",		-- 8, 9, 9, 9
        5370 => x"09000000",		-- 9, 8, 8, 8
        5371 => x"00000000",		-- 8, 8, 8, 8
        5372 => x"00000009",		-- 8, 8, 8, 9
        5373 => x"09090909",		-- 9, 9, 9, 9
        5374 => x"0B0B0B0B",		-- 11, 11, 11, 11
        5375 => x"00000000",		-- 8, 8, 8, 8
        5376 => x"00090909",		-- 8, 9, 9, 9
        5377 => x"0A09090B",		-- 10, 9, 9, 11
        5378 => x"0B0B0B0B",		-- 11, 11, 11, 11
        5379 => x"0B000000",		-- 11, 8, 8, 8
        5380 => x"09090909",		-- 9, 9, 9, 9
        5381 => x"0A0A0B0B",		-- 10, 10, 11, 11
        5382 => x"0B0B0B0B",		-- 11, 11, 11, 11
        5383 => x"00000000",		-- 8, 8, 8, 8
        5384 => x"09000909",		-- 9, 8, 9, 9
        5385 => x"0A0A0A0B",		-- 10, 10, 10, 11
        5386 => x"0A0A090A",		-- 10, 10, 9, 10
        5387 => x"00000000",		-- 8, 8, 8, 8
        5388 => x"0000090B",		-- 8, 8, 9, 11
        5389 => x"0B0A0A0B",		-- 11, 10, 10, 11
        5390 => x"0A0A0B0A",		-- 10, 10, 11, 10
        5391 => x"0A0A0000",		-- 10, 10, 8, 8
        5392 => x"0000000B",		-- 8, 8, 8, 11
        5393 => x"0B0B0A0A",		-- 11, 11, 10, 10
        5394 => x"0A0A0A0A",		-- 10, 10, 10, 10
        5395 => x"000B0000",		-- 8, 11, 8, 8
        5396 => x"00000000",		-- 8, 8, 8, 8
        5397 => x"09090909",		-- 9, 9, 9, 9
        5398 => x"0A0A0A0A",		-- 10, 10, 10, 10
        5399 => x"000B0000",		-- 8, 11, 8, 8
        5400 => x"0000090B",		-- 8, 8, 9, 11
        5401 => x"0B09090A",		-- 11, 9, 9, 10
        5402 => x"0A0A0B0B",		-- 10, 10, 11, 11
        5403 => x"0A0B0000",		-- 10, 11, 8, 8
        5404 => x"00000B0B",		-- 8, 8, 11, 11
        5405 => x"0B0B0B0A",		-- 11, 11, 11, 10
        5406 => x"0A0A090B",		-- 10, 10, 9, 11
        5407 => x"0A0B0000",		-- 10, 11, 8, 8
        5408 => x"00090B0B",		-- 8, 9, 11, 11
        5409 => x"0B0B0B0A",		-- 11, 11, 11, 10
        5410 => x"0A09090B",		-- 10, 9, 9, 11
        5411 => x"000B0000",		-- 8, 11, 8, 8
        5412 => x"0009090B",		-- 8, 9, 9, 11
        5413 => x"0B0B0B09",		-- 11, 11, 11, 9
        5414 => x"09090B00",		-- 9, 9, 11, 8
        5415 => x"000B0000",		-- 8, 11, 8, 8
        5416 => x"0B0B0909",		-- 11, 11, 9, 9
        5417 => x"0909090B",		-- 9, 9, 9, 11
        5418 => x"0B0B0B09",		-- 11, 11, 11, 9
        5419 => x"000B0000",		-- 8, 11, 8, 8
        5420 => x"0B0B0B09",		-- 11, 11, 11, 9
        5421 => x"09090909",		-- 9, 9, 9, 9
        5422 => x"0909090B",		-- 9, 9, 9, 11
        5423 => x"0B000000",		-- 11, 8, 8, 8
        5424 => x"000B0B0B",		-- 8, 11, 11, 11
        5425 => x"00000000",		-- 8, 8, 8, 8
        5426 => x"000B0B0B",		-- 8, 11, 11, 11
        5427 => x"00000000",		-- 8, 8, 8, 8

                --  sprite 4
        5428 => x"00000000",		-- 8, 8, 8, 8
        5429 => x"00090909",		-- 8, 9, 9, 9
        5430 => x"09000000",		-- 9, 8, 8, 8
        5431 => x"00000000",		-- 8, 8, 8, 8
        5432 => x"00000009",		-- 8, 8, 8, 9
        5433 => x"09090909",		-- 9, 9, 9, 9
        5434 => x"0B0B0B0B",		-- 11, 11, 11, 11
        5435 => x"00000000",		-- 8, 8, 8, 8
        5436 => x"00090909",		-- 8, 9, 9, 9
        5437 => x"0A09090B",		-- 10, 9, 9, 11
        5438 => x"0B0B0B0B",		-- 11, 11, 11, 11
        5439 => x"0B000000",		-- 11, 8, 8, 8
        5440 => x"09090909",		-- 9, 9, 9, 9
        5441 => x"0A0A0B0B",		-- 10, 10, 11, 11
        5442 => x"0B0B0B0B",		-- 11, 11, 11, 11
        5443 => x"00000000",		-- 8, 8, 8, 8
        5444 => x"09000909",		-- 9, 8, 9, 9
        5445 => x"0A0A0A0B",		-- 10, 10, 10, 11
        5446 => x"0A0A090A",		-- 10, 10, 9, 10
        5447 => x"00000B00",		-- 8, 8, 11, 8
        5448 => x"0000090B",		-- 8, 8, 9, 11
        5449 => x"0B0A0A0B",		-- 11, 10, 10, 11
        5450 => x"0A0A0B0A",		-- 10, 10, 11, 10
        5451 => x"0A0A0B00",		-- 10, 10, 11, 8
        5452 => x"0000000B",		-- 8, 8, 8, 11
        5453 => x"0B0B0A0A",		-- 11, 11, 10, 10
        5454 => x"0A0A0A0A",		-- 10, 10, 10, 10
        5455 => x"00000B00",		-- 8, 8, 11, 8
        5456 => x"00000000",		-- 8, 8, 8, 8
        5457 => x"09090909",		-- 9, 9, 9, 9
        5458 => x"0A0A0A0A",		-- 10, 10, 10, 10
        5459 => x"00000B00",		-- 8, 8, 11, 8
        5460 => x"00000B09",		-- 8, 8, 11, 9
        5461 => x"09090909",		-- 9, 9, 9, 9
        5462 => x"09090B0B",		-- 9, 9, 11, 11
        5463 => x"0B0A0B00",		-- 11, 10, 11, 8
        5464 => x"000B0B0B",		-- 8, 11, 11, 11
        5465 => x"090A0A0A",		-- 9, 10, 10, 10
        5466 => x"0909090B",		-- 9, 9, 9, 11
        5467 => x"0B0A0B00",		-- 11, 10, 11, 8
        5468 => x"000B0B0B",		-- 8, 11, 11, 11
        5469 => x"0B0A0A0A",		-- 11, 10, 10, 10
        5470 => x"0909090B",		-- 9, 9, 9, 11
        5471 => x"0B000B00",		-- 11, 8, 11, 8
        5472 => x"000B0B0B",		-- 8, 11, 11, 11
        5473 => x"0B0A0A09",		-- 11, 10, 10, 9
        5474 => x"09090B00",		-- 9, 9, 11, 8
        5475 => x"00000B00",		-- 8, 8, 11, 8
        5476 => x"0000090B",		-- 8, 8, 9, 11
        5477 => x"0B09090B",		-- 11, 9, 9, 11
        5478 => x"0B0B0B00",		-- 11, 11, 11, 8
        5479 => x"00000B00",		-- 8, 8, 11, 8
        5480 => x"00090909",		-- 8, 9, 9, 9
        5481 => x"09090909",		-- 9, 9, 9, 9
        5482 => x"09090900",		-- 9, 9, 9, 8
        5483 => x"00000000",		-- 8, 8, 8, 8
        5484 => x"00000000",		-- 8, 8, 8, 8
        5485 => x"0B0B0B0B",		-- 11, 11, 11, 11
        5486 => x"00000000",		-- 8, 8, 8, 8
        5487 => x"00000000",		-- 8, 8, 8, 8
        5488 => x"00000000",		-- 8, 8, 8, 8
        5489 => x"0B0B0B0B",		-- 11, 11, 11, 11
        5490 => x"0B000000",		-- 11, 8, 8, 8
        5491 => x"00000000",		-- 8, 8, 8, 8

                --  sprite 5
        5492 => x"00000000",		-- 8, 8, 8, 8
        5493 => x"00090909",		-- 8, 9, 9, 9
        5494 => x"09090900",		-- 9, 9, 9, 8
        5495 => x"00000000",		-- 8, 8, 8, 8
        5496 => x"00000000",		-- 8, 8, 8, 8
        5497 => x"09090909",		-- 9, 9, 9, 9
        5498 => x"09090909",		-- 9, 9, 9, 9
        5499 => x"00000000",		-- 8, 8, 8, 8
        5500 => x"00000A00",		-- 8, 8, 10, 8
        5501 => x"090B0B0B",		-- 9, 11, 11, 11
        5502 => x"0B0B0B09",		-- 11, 11, 11, 9
        5503 => x"000A0000",		-- 8, 10, 8, 8
        5504 => x"00000A00",		-- 8, 8, 10, 8
        5505 => x"0B0B0B0B",		-- 11, 11, 11, 11
        5506 => x"0B0B0B0B",		-- 11, 11, 11, 11
        5507 => x"000A0000",		-- 8, 10, 8, 8
        5508 => x"00000A0A",		-- 8, 8, 10, 10
        5509 => x"0B0A090A",		-- 11, 10, 9, 10
        5510 => x"0A090A0B",		-- 10, 9, 10, 11
        5511 => x"0A0A0000",		-- 10, 10, 8, 8
        5512 => x"00000A0A",		-- 8, 8, 10, 10
        5513 => x"0B0A0B0A",		-- 11, 10, 11, 10
        5514 => x"0A0B0A0B",		-- 10, 11, 10, 11
        5515 => x"0A0A0000",		-- 10, 10, 8, 8
        5516 => x"0B0B0B0B",		-- 11, 11, 11, 11
        5517 => x"0B0B0B0B",		-- 11, 11, 11, 11
        5518 => x"0A0A0A0A",		-- 10, 10, 10, 10
        5519 => x"0A0B0000",		-- 10, 11, 8, 8
        5520 => x"0B0B0B0A",		-- 11, 11, 11, 10
        5521 => x"0A0B0B0B",		-- 10, 11, 11, 11
        5522 => x"0B0A0A09",		-- 11, 10, 10, 9
        5523 => x"090B0000",		-- 9, 11, 8, 8
        5524 => x"0B0B0B0A",		-- 11, 11, 11, 10
        5525 => x"0A0B0B0B",		-- 10, 11, 11, 11
        5526 => x"0A0A0909",		-- 10, 10, 9, 9
        5527 => x"0B0B0B00",		-- 11, 11, 11, 8
        5528 => x"0B0A0A0A",		-- 11, 10, 10, 10
        5529 => x"0A0A0A0B",		-- 10, 10, 10, 11
        5530 => x"09090909",		-- 9, 9, 9, 9
        5531 => x"0A0B0B00",		-- 10, 11, 11, 8
        5532 => x"0B0A0A0A",		-- 11, 10, 10, 10
        5533 => x"0A0A0A0B",		-- 10, 10, 10, 11
        5534 => x"0B09090A",		-- 11, 9, 9, 10
        5535 => x"0A0A0B00",		-- 10, 10, 11, 8
        5536 => x"0B0B0B0A",		-- 11, 11, 11, 10
        5537 => x"0A0B0B0B",		-- 10, 11, 11, 11
        5538 => x"0B0B0B0B",		-- 11, 11, 11, 11
        5539 => x"0A0A0A00",		-- 10, 10, 10, 8
        5540 => x"0B0B0B0A",		-- 11, 11, 11, 10
        5541 => x"0A0B0B0B",		-- 10, 11, 11, 11
        5542 => x"0B090909",		-- 11, 9, 9, 9
        5543 => x"090A0000",		-- 9, 10, 8, 8
        5544 => x"0B0B0B0A",		-- 11, 11, 11, 10
        5545 => x"0A0B0B0B",		-- 10, 11, 11, 11
        5546 => x"09090909",		-- 9, 9, 9, 9
        5547 => x"00000000",		-- 8, 8, 8, 8
        5548 => x"000B0B0B",		-- 8, 11, 11, 11
        5549 => x"0B0B0B00",		-- 11, 11, 11, 8
        5550 => x"000B0B0B",		-- 8, 11, 11, 11
        5551 => x"00000000",		-- 8, 8, 8, 8
        5552 => x"00000B0B",		-- 8, 8, 11, 11
        5553 => x"0B0B0000",		-- 11, 11, 8, 8
        5554 => x"00000000",		-- 8, 8, 8, 8
        5555 => x"00000000",		-- 8, 8, 8, 8

                --  sprite 6
        5556 => x"00000000",		-- 8, 8, 8, 8
        5557 => x"00090909",		-- 8, 9, 9, 9
        5558 => x"09090900",		-- 9, 9, 9, 8
        5559 => x"00000000",		-- 8, 8, 8, 8
        5560 => x"00000000",		-- 8, 8, 8, 8
        5561 => x"09090909",		-- 9, 9, 9, 9
        5562 => x"09090909",		-- 9, 9, 9, 9
        5563 => x"00000000",		-- 8, 8, 8, 8
        5564 => x"00000A00",		-- 8, 8, 10, 8
        5565 => x"090B0B0B",		-- 9, 11, 11, 11
        5566 => x"0B0B0B09",		-- 11, 11, 11, 9
        5567 => x"000A0000",		-- 8, 10, 8, 8
        5568 => x"00000A00",		-- 8, 8, 10, 8
        5569 => x"0B0B0B0B",		-- 11, 11, 11, 11
        5570 => x"0B0B0B0B",		-- 11, 11, 11, 11
        5571 => x"000A0000",		-- 8, 10, 8, 8
        5572 => x"00000A0A",		-- 8, 8, 10, 10
        5573 => x"0B0A090A",		-- 11, 10, 9, 10
        5574 => x"0A090A0B",		-- 10, 9, 10, 11
        5575 => x"0A0A0000",		-- 10, 10, 8, 8
        5576 => x"00000A0A",		-- 8, 8, 10, 10
        5577 => x"0B0A0B0A",		-- 11, 10, 11, 10
        5578 => x"0A0B0A0B",		-- 10, 11, 10, 11
        5579 => x"0A0A0000",		-- 10, 10, 8, 8
        5580 => x"0B0B0B0B",		-- 11, 11, 11, 11
        5581 => x"0B0B0B0B",		-- 11, 11, 11, 11
        5582 => x"0A0A0A0A",		-- 10, 10, 10, 10
        5583 => x"0A0B0000",		-- 10, 11, 8, 8
        5584 => x"0B0B0B0A",		-- 11, 11, 11, 10
        5585 => x"0A0B0B0B",		-- 10, 11, 11, 11
        5586 => x"0B0A0A09",		-- 11, 10, 10, 9
        5587 => x"0B0B0000",		-- 11, 11, 8, 8
        5588 => x"0B0B0B0A",		-- 11, 11, 11, 10
        5589 => x"0A0B0B0B",		-- 10, 11, 11, 11
        5590 => x"0A0A0909",		-- 10, 10, 9, 9
        5591 => x"090A0000",		-- 9, 10, 8, 8
        5592 => x"0B0A0A0A",		-- 11, 10, 10, 10
        5593 => x"0A0A0A0B",		-- 10, 10, 10, 11
        5594 => x"09090909",		-- 9, 9, 9, 9
        5595 => x"090A0000",		-- 9, 10, 8, 8
        5596 => x"0B0A0A0A",		-- 11, 10, 10, 10
        5597 => x"0A0A0A0B",		-- 10, 10, 10, 11
        5598 => x"0B0B0909",		-- 11, 11, 9, 9
        5599 => x"0B000000",		-- 11, 8, 8, 8
        5600 => x"0B0B0B0A",		-- 11, 11, 11, 10
        5601 => x"0A0B0B0B",		-- 10, 11, 11, 11
        5602 => x"090B0B0B",		-- 9, 11, 11, 11
        5603 => x"09000000",		-- 9, 8, 8, 8
        5604 => x"0B0B0B0A",		-- 11, 11, 11, 10
        5605 => x"0A0B0B0B",		-- 10, 11, 11, 11
        5606 => x"0B0B0909",		-- 11, 11, 9, 9
        5607 => x"09000000",		-- 9, 8, 8, 8
        5608 => x"0B0B0B0A",		-- 11, 11, 11, 10
        5609 => x"0A0B0B0B",		-- 10, 11, 11, 11
        5610 => x"0909090B",		-- 9, 9, 9, 11
        5611 => x"00000000",		-- 8, 8, 8, 8
        5612 => x"000B0B0B",		-- 8, 11, 11, 11
        5613 => x"0B0B0B00",		-- 11, 11, 11, 8
        5614 => x"000B0B0B",		-- 8, 11, 11, 11
        5615 => x"00000000",		-- 8, 8, 8, 8
        5616 => x"00000B0B",		-- 8, 8, 11, 11
        5617 => x"0B0B0000",		-- 11, 11, 8, 8
        5618 => x"000B0B0B",		-- 8, 11, 11, 11
        5619 => x"00000000",		-- 8, 8, 8, 8

                --  sprite 7
        5620 => x"00000000",		-- 8, 8, 8, 8
        5621 => x"00000000",		-- 8, 8, 8, 8
        5622 => x"00000000",		-- 8, 8, 8, 8
        5623 => x"00000000",		-- 8, 8, 8, 8
        5624 => x"00000000",		-- 8, 8, 8, 8
        5625 => x"00090909",		-- 8, 9, 9, 9
        5626 => x"09000000",		-- 9, 8, 8, 8
        5627 => x"00000000",		-- 8, 8, 8, 8
        5628 => x"00000009",		-- 8, 8, 8, 9
        5629 => x"09090909",		-- 9, 9, 9, 9
        5630 => x"0B0B0B0B",		-- 11, 11, 11, 11
        5631 => x"00000000",		-- 8, 8, 8, 8
        5632 => x"00090909",		-- 8, 9, 9, 9
        5633 => x"0A09090B",		-- 10, 9, 9, 11
        5634 => x"0B0B0B0B",		-- 11, 11, 11, 11
        5635 => x"0B000000",		-- 11, 8, 8, 8
        5636 => x"09090909",		-- 9, 9, 9, 9
        5637 => x"0A0A0B0B",		-- 10, 10, 11, 11
        5638 => x"0B0B0B0B",		-- 11, 11, 11, 11
        5639 => x"000B0B00",		-- 8, 11, 11, 8
        5640 => x"09000909",		-- 9, 8, 9, 9
        5641 => x"0A0A0A0B",		-- 10, 10, 10, 11
        5642 => x"0A0A090A",		-- 10, 10, 9, 10
        5643 => x"000B0B00",		-- 8, 11, 11, 8
        5644 => x"0000090B",		-- 8, 8, 9, 11
        5645 => x"0B0A0A0B",		-- 11, 10, 10, 11
        5646 => x"0A0A0B0A",		-- 10, 10, 11, 10
        5647 => x"0A0B0A00",		-- 10, 11, 10, 8
        5648 => x"0000000B",		-- 8, 8, 8, 11
        5649 => x"0B0B0A0A",		-- 11, 11, 10, 10
        5650 => x"0A0A0A0A",		-- 10, 10, 10, 10
        5651 => x"000B0A00",		-- 8, 11, 10, 8
        5652 => x"00000000",		-- 8, 8, 8, 8
        5653 => x"09090909",		-- 9, 9, 9, 9
        5654 => x"0A0A0A0A",		-- 10, 10, 10, 10
        5655 => x"000B0A00",		-- 8, 11, 10, 8
        5656 => x"0000090B",		-- 8, 8, 9, 11
        5657 => x"0B09090A",		-- 11, 9, 9, 10
        5658 => x"0A0A0B0B",		-- 10, 10, 11, 11
        5659 => x"0A0B0A00",		-- 10, 11, 10, 8
        5660 => x"00000B0B",		-- 8, 8, 11, 11
        5661 => x"0B0B0B0A",		-- 11, 11, 11, 10
        5662 => x"0A0A090B",		-- 10, 10, 9, 11
        5663 => x"0A0B0A00",		-- 10, 11, 10, 8
        5664 => x"00090B0B",		-- 8, 9, 11, 11
        5665 => x"0B0B0B0A",		-- 11, 11, 11, 10
        5666 => x"0A09090B",		-- 10, 9, 9, 11
        5667 => x"000B0A00",		-- 8, 11, 10, 8
        5668 => x"0009090B",		-- 8, 9, 9, 11
        5669 => x"0B0B0B09",		-- 11, 11, 11, 9
        5670 => x"09090B00",		-- 9, 9, 11, 8
        5671 => x"000B0A00",		-- 8, 11, 10, 8
        5672 => x"0B0B0909",		-- 11, 11, 9, 9
        5673 => x"0909090B",		-- 9, 9, 9, 11
        5674 => x"0B0B0B09",		-- 11, 11, 11, 9
        5675 => x"000B0A00",		-- 8, 11, 10, 8
        5676 => x"0B0B0B09",		-- 11, 11, 11, 9
        5677 => x"09090909",		-- 9, 9, 9, 9
        5678 => x"0909090B",		-- 9, 9, 9, 11
        5679 => x"0B0B0B00",		-- 11, 11, 11, 8
        5680 => x"000B0B0B",		-- 8, 11, 11, 11
        5681 => x"00000000",		-- 8, 8, 8, 8
        5682 => x"000B0B0B",		-- 8, 11, 11, 11
        5683 => x"000B0B00",		-- 8, 11, 11, 8

                --  sprite 8
        5684 => x"00000000",		-- 8, 8, 8, 8
        5685 => x"00090909",		-- 8, 9, 9, 9
        5686 => x"09000000",		-- 9, 8, 8, 8
        5687 => x"00000000",		-- 8, 8, 8, 8
        5688 => x"00000009",		-- 8, 8, 8, 9
        5689 => x"09090909",		-- 9, 9, 9, 9
        5690 => x"0B0B0B0B",		-- 11, 11, 11, 11
        5691 => x"00000000",		-- 8, 8, 8, 8
        5692 => x"00090909",		-- 8, 9, 9, 9
        5693 => x"0A09090B",		-- 10, 9, 9, 11
        5694 => x"0B0B0B0B",		-- 11, 11, 11, 11
        5695 => x"0B000000",		-- 11, 8, 8, 8
        5696 => x"09090909",		-- 9, 9, 9, 9
        5697 => x"0A0A0B0B",		-- 10, 10, 11, 11
        5698 => x"0B0B0B0B",		-- 11, 11, 11, 11
        5699 => x"00000B0B",		-- 8, 8, 11, 11
        5700 => x"09000909",		-- 9, 8, 9, 9
        5701 => x"0A0A0A0B",		-- 10, 10, 10, 11
        5702 => x"0A0A090A",		-- 10, 10, 9, 10
        5703 => x"00000B0B",		-- 8, 8, 11, 11
        5704 => x"0000090B",		-- 8, 8, 9, 11
        5705 => x"0B0A0A0B",		-- 11, 10, 10, 11
        5706 => x"0A0A0B0A",		-- 10, 10, 11, 10
        5707 => x"0A0A0B0A",		-- 10, 10, 11, 10
        5708 => x"0000000B",		-- 8, 8, 8, 11
        5709 => x"0B0B0A0A",		-- 11, 11, 10, 10
        5710 => x"0A0A0A0A",		-- 10, 10, 10, 10
        5711 => x"00000B0A",		-- 8, 8, 11, 10
        5712 => x"00000000",		-- 8, 8, 8, 8
        5713 => x"09090909",		-- 9, 9, 9, 9
        5714 => x"0A0A0A0A",		-- 10, 10, 10, 10
        5715 => x"00000B0A",		-- 8, 8, 11, 10
        5716 => x"00000B09",		-- 8, 8, 11, 9
        5717 => x"09090909",		-- 9, 9, 9, 9
        5718 => x"09090B0B",		-- 9, 9, 11, 11
        5719 => x"0B0A0B0A",		-- 11, 10, 11, 10
        5720 => x"000B0B0B",		-- 8, 11, 11, 11
        5721 => x"090A0A0A",		-- 9, 10, 10, 10
        5722 => x"0909090B",		-- 9, 9, 9, 11
        5723 => x"0B0A0B0A",		-- 11, 10, 11, 10
        5724 => x"000B0B0B",		-- 8, 11, 11, 11
        5725 => x"0B0A0A0A",		-- 11, 10, 10, 10
        5726 => x"0909090B",		-- 9, 9, 9, 11
        5727 => x"0B000B0A",		-- 11, 8, 11, 10
        5728 => x"000B0B0B",		-- 8, 11, 11, 11
        5729 => x"0B0A0A09",		-- 11, 10, 10, 9
        5730 => x"09090B00",		-- 9, 9, 11, 8
        5731 => x"00000B0A",		-- 8, 8, 11, 10
        5732 => x"0000090B",		-- 8, 8, 9, 11
        5733 => x"0B09090B",		-- 11, 9, 9, 11
        5734 => x"0B0B0B00",		-- 11, 11, 11, 8
        5735 => x"00000B0A",		-- 8, 8, 11, 10
        5736 => x"00090909",		-- 8, 9, 9, 9
        5737 => x"09090909",		-- 9, 9, 9, 9
        5738 => x"09090900",		-- 9, 9, 9, 8
        5739 => x"00000B0B",		-- 8, 8, 11, 11
        5740 => x"00000000",		-- 8, 8, 8, 8
        5741 => x"0B0B0B0B",		-- 11, 11, 11, 11
        5742 => x"00000000",		-- 8, 8, 8, 8
        5743 => x"00000B0B",		-- 8, 8, 11, 11
        5744 => x"00000000",		-- 8, 8, 8, 8
        5745 => x"0B0B0B0B",		-- 11, 11, 11, 11
        5746 => x"0B000000",		-- 11, 8, 8, 8
        5747 => x"00000000",		-- 8, 8, 8, 8

                --  sprite 9
        5748 => x"0000000B",		-- 8, 8, 8, 11
        5749 => x"0B000909",		-- 11, 8, 9, 9
        5750 => x"09090900",		-- 9, 9, 9, 8
        5751 => x"00000000",		-- 8, 8, 8, 8
        5752 => x"00000B0A",		-- 8, 8, 11, 10
        5753 => x"0B090909",		-- 11, 9, 9, 9
        5754 => x"09090909",		-- 9, 9, 9, 9
        5755 => x"00000000",		-- 8, 8, 8, 8
        5756 => x"000B0B0A",		-- 8, 11, 11, 10
        5757 => x"09090B0B",		-- 9, 9, 11, 11
        5758 => x"0B0B0909",		-- 11, 11, 9, 9
        5759 => x"09000000",		-- 9, 8, 8, 8
        5760 => x"0B0B0A0A",		-- 11, 11, 10, 10
        5761 => x"090B0B0B",		-- 9, 11, 11, 11
        5762 => x"0B0B0B09",		-- 11, 11, 11, 9
        5763 => x"09000A00",		-- 9, 8, 10, 8
        5764 => x"0B0B0A0A",		-- 11, 11, 10, 10
        5765 => x"0B0A090A",		-- 11, 10, 9, 10
        5766 => x"0A090B0B",		-- 10, 9, 11, 11
        5767 => x"090A0A00",		-- 9, 10, 10, 8
        5768 => x"0A0B0B0A",		-- 10, 11, 11, 10
        5769 => x"0B0A0B0A",		-- 11, 10, 11, 10
        5770 => x"0A0B0A0B",		-- 10, 11, 10, 11
        5771 => x"090A0000",		-- 9, 10, 8, 8
        5772 => x"000A0B0B",		-- 8, 10, 11, 11
        5773 => x"090A0A0B",		-- 9, 10, 10, 11
        5774 => x"0B0A0A0A",		-- 11, 10, 10, 10
        5775 => x"0A000000",		-- 10, 8, 8, 8
        5776 => x"00000A0B",		-- 8, 8, 10, 11
        5777 => x"09090A0B",		-- 9, 9, 10, 11
        5778 => x"0B0A0A0B",		-- 11, 10, 10, 11
        5779 => x"0B000000",		-- 11, 8, 8, 8
        5780 => x"0000000A",		-- 8, 8, 8, 10
        5781 => x"0909090A",		-- 9, 9, 9, 10
        5782 => x"0A0A0B0B",		-- 10, 10, 11, 11
        5783 => x"0B0B0000",		-- 11, 11, 8, 8
        5784 => x"00000000",		-- 8, 8, 8, 8
        5785 => x"0B090909",		-- 11, 9, 9, 9
        5786 => x"09090B0B",		-- 9, 9, 11, 11
        5787 => x"0B0B0000",		-- 11, 11, 8, 8
        5788 => x"00000000",		-- 8, 8, 8, 8
        5789 => x"090B090B",		-- 9, 11, 9, 11
        5790 => x"0B0B0B0B",		-- 11, 11, 11, 11
        5791 => x"0B090000",		-- 11, 9, 8, 8
        5792 => x"00000000",		-- 8, 8, 8, 8
        5793 => x"09090B0B",		-- 9, 9, 11, 11
        5794 => x"090B0B0B",		-- 9, 11, 11, 11
        5795 => x"09090000",		-- 9, 9, 8, 8
        5796 => x"0000000B",		-- 8, 8, 8, 11
        5797 => x"0B09090B",		-- 11, 9, 9, 11
        5798 => x"0B0A0A0B",		-- 11, 10, 10, 11
        5799 => x"09090B00",		-- 9, 9, 11, 8
        5800 => x"00000B0B",		-- 8, 8, 11, 11
        5801 => x"0B000909",		-- 11, 8, 9, 9
        5802 => x"0A0A0A09",		-- 10, 10, 10, 9
        5803 => x"090B0B0B",		-- 9, 11, 11, 11
        5804 => x"00000000",		-- 8, 8, 8, 8
        5805 => x"00000000",		-- 8, 8, 8, 8
        5806 => x"0A0A0A00",		-- 10, 10, 10, 8
        5807 => x"0B0B0B0B",		-- 11, 11, 11, 11
        5808 => x"00000000",		-- 8, 8, 8, 8
        5809 => x"00000000",		-- 8, 8, 8, 8
        5810 => x"00000000",		-- 8, 8, 8, 8
        5811 => x"00000000",		-- 8, 8, 8, 8

                --  sprite 10
        5812 => x"0000000B",		-- 8, 8, 8, 11
        5813 => x"09090909",		-- 9, 9, 9, 9
        5814 => x"09000000",		-- 9, 8, 8, 8
        5815 => x"00000000",		-- 8, 8, 8, 8
        5816 => x"000A0009",		-- 8, 10, 8, 9
        5817 => x"09090909",		-- 9, 9, 9, 9
        5818 => x"09090000",		-- 9, 9, 8, 8
        5819 => x"00000000",		-- 8, 8, 8, 8
        5820 => x"000A0B09",		-- 8, 10, 11, 9
        5821 => x"09090909",		-- 9, 9, 9, 9
        5822 => x"09090900",		-- 9, 9, 9, 8
        5823 => x"00000000",		-- 8, 8, 8, 8
        5824 => x"000A0A09",		-- 8, 10, 10, 9
        5825 => x"09090909",		-- 9, 9, 9, 9
        5826 => x"09090900",		-- 9, 9, 9, 8
        5827 => x"0A000000",		-- 10, 8, 8, 8
        5828 => x"000B0A0B",		-- 8, 11, 10, 11
        5829 => x"09090909",		-- 9, 9, 9, 9
        5830 => x"09090B0A",		-- 9, 9, 11, 10
        5831 => x"0A000000",		-- 10, 8, 8, 8
        5832 => x"000B0A0B",		-- 8, 11, 10, 11
        5833 => x"0B090909",		-- 11, 9, 9, 9
        5834 => x"0B0B0B0A",		-- 11, 11, 11, 10
        5835 => x"0000000A",		-- 8, 8, 8, 10
        5836 => x"000B0B09",		-- 8, 11, 11, 9
        5837 => x"0B0B090B",		-- 11, 11, 9, 11
        5838 => x"0B0B090A",		-- 11, 11, 9, 10
        5839 => x"00000A0B",		-- 8, 8, 10, 11
        5840 => x"000B0B09",		-- 8, 11, 11, 9
        5841 => x"090B0B0B",		-- 9, 11, 11, 11
        5842 => x"0B090B0B",		-- 11, 9, 11, 11
        5843 => x"0B0A0B0B",		-- 11, 10, 11, 11
        5844 => x"00000B09",		-- 8, 8, 11, 9
        5845 => x"09090909",		-- 9, 9, 9, 9
        5846 => x"09090B0B",		-- 9, 9, 11, 11
        5847 => x"0A0B0B0B",		-- 10, 11, 11, 11
        5848 => x"00000B09",		-- 8, 8, 11, 9
        5849 => x"09090909",		-- 9, 9, 9, 9
        5850 => x"09090B0A",		-- 9, 9, 11, 10
        5851 => x"0B0B0B0B",		-- 11, 11, 11, 11
        5852 => x"0000090B",		-- 8, 8, 9, 11
        5853 => x"09090909",		-- 9, 9, 9, 9
        5854 => x"09090A0B",		-- 9, 9, 10, 11
        5855 => x"0B0B0B00",		-- 11, 11, 11, 8
        5856 => x"000B0909",		-- 8, 11, 9, 9
        5857 => x"0B0B0B0B",		-- 11, 11, 11, 11
        5858 => x"0B0B0B0A",		-- 11, 11, 11, 10
        5859 => x"0B0B0000",		-- 11, 11, 8, 8
        5860 => x"0B0B0909",		-- 11, 11, 9, 9
        5861 => x"09090909",		-- 9, 9, 9, 9
        5862 => x"09090909",		-- 9, 9, 9, 9
        5863 => x"0A000000",		-- 10, 8, 8, 8
        5864 => x"0B0B0B00",		-- 11, 11, 11, 8
        5865 => x"00000009",		-- 8, 8, 8, 9
        5866 => x"0909090B",		-- 9, 9, 9, 11
        5867 => x"0B000000",		-- 11, 8, 8, 8
        5868 => x"00000000",		-- 8, 8, 8, 8
        5869 => x"00000000",		-- 8, 8, 8, 8
        5870 => x"00000B0B",		-- 8, 8, 11, 11
        5871 => x"0B0B0000",		-- 11, 11, 8, 8
        5872 => x"00000000",		-- 8, 8, 8, 8
        5873 => x"00000000",		-- 8, 8, 8, 8
        5874 => x"00000B0B",		-- 8, 8, 11, 11
        5875 => x"0B0B0000",		-- 11, 11, 8, 8

                --  sprite 11
        5876 => x"00000000",		-- 8, 8, 8, 8
        5877 => x"00000000",		-- 8, 8, 8, 8
        5878 => x"00000000",		-- 8, 8, 8, 8
        5879 => x"00000000",		-- 8, 8, 8, 8
        5880 => x"00000000",		-- 8, 8, 8, 8
        5881 => x"00000909",		-- 8, 8, 9, 9
        5882 => x"09090000",		-- 9, 9, 8, 8
        5883 => x"00000000",		-- 8, 8, 8, 8
        5884 => x"00000000",		-- 8, 8, 8, 8
        5885 => x"09090909",		-- 9, 9, 9, 9
        5886 => x"090B0B0B",		-- 9, 11, 11, 11
        5887 => x"0B000000",		-- 11, 8, 8, 8
        5888 => x"00000009",		-- 8, 8, 8, 9
        5889 => x"090A0909",		-- 9, 10, 9, 9
        5890 => x"0B0B0B0B",		-- 11, 11, 11, 11
        5891 => x"0B0B0000",		-- 11, 11, 8, 8
        5892 => x"00000009",		-- 8, 8, 8, 9
        5893 => x"090A0A0B",		-- 9, 10, 10, 11
        5894 => x"0B0B0B0B",		-- 11, 11, 11, 11
        5895 => x"0B000000",		-- 11, 8, 8, 8
        5896 => x"00000909",		-- 8, 8, 9, 9
        5897 => x"090A0A0A",		-- 9, 10, 10, 10
        5898 => x"0B0A0A09",		-- 11, 10, 10, 9
        5899 => x"0A000000",		-- 10, 8, 8, 8
        5900 => x"00090909",		-- 8, 9, 9, 9
        5901 => x"0B0B0A0A",		-- 11, 11, 10, 10
        5902 => x"0B0A0A0B",		-- 11, 10, 10, 11
        5903 => x"0A0A0A00",		-- 10, 10, 10, 8
        5904 => x"00090000",		-- 8, 9, 8, 8
        5905 => x"0B0B0B0A",		-- 11, 11, 11, 10
        5906 => x"0A0A0A0A",		-- 10, 10, 10, 10
        5907 => x"0A000000",		-- 10, 8, 8, 8
        5908 => x"00000000",		-- 8, 8, 8, 8
        5909 => x"09090909",		-- 9, 9, 9, 9
        5910 => x"090A0A0A",		-- 9, 10, 10, 10
        5911 => x"0A0A0000",		-- 10, 10, 8, 8
        5912 => x"00000009",		-- 8, 8, 8, 9
        5913 => x"090B0B0B",		-- 9, 11, 11, 11
        5914 => x"0B0B0B0A",		-- 11, 11, 11, 10
        5915 => x"0A0A0000",		-- 10, 10, 8, 8
        5916 => x"00000009",		-- 8, 8, 8, 9
        5917 => x"0B0B0B0B",		-- 11, 11, 11, 11
        5918 => x"0B0B0B0A",		-- 11, 11, 11, 10
        5919 => x"0A000000",		-- 10, 8, 8, 8
        5920 => x"00000909",		-- 8, 8, 9, 9
        5921 => x"0B0B0B0B",		-- 11, 11, 11, 11
        5922 => x"0B0B0B09",		-- 11, 11, 11, 9
        5923 => x"00000000",		-- 8, 8, 8, 8
        5924 => x"00090909",		-- 8, 9, 9, 9
        5925 => x"090B0B0B",		-- 9, 11, 11, 11
        5926 => x"0909090B",		-- 9, 9, 9, 11
        5927 => x"0B000000",		-- 11, 8, 8, 8
        5928 => x"0B0B0909",		-- 11, 11, 9, 9
        5929 => x"09090909",		-- 9, 9, 9, 9
        5930 => x"0B0B0B0B",		-- 11, 11, 11, 11
        5931 => x"0B000000",		-- 11, 8, 8, 8
        5932 => x"0B0B0B09",		-- 11, 11, 11, 9
        5933 => x"09090909",		-- 9, 9, 9, 9
        5934 => x"09090909",		-- 9, 9, 9, 9
        5935 => x"0B0B0000",		-- 11, 11, 8, 8
        5936 => x"000B0B0B",		-- 8, 11, 11, 11
        5937 => x"00000000",		-- 8, 8, 8, 8
        5938 => x"0000000B",		-- 8, 8, 8, 11
        5939 => x"0B0B0B00",		-- 11, 11, 11, 8

                --  sprite 12
        5940 => x"000A0A00",		-- 8, 10, 10, 8
        5941 => x"00000909",		-- 8, 8, 9, 9
        5942 => x"09090900",		-- 9, 9, 9, 8
        5943 => x"00000000",		-- 8, 8, 8, 8
        5944 => x"000A0A0A",		-- 8, 10, 10, 10
        5945 => x"00090B0B",		-- 8, 9, 11, 11
        5946 => x"09090909",		-- 9, 9, 9, 9
        5947 => x"00000000",		-- 8, 8, 8, 8
        5948 => x"000B0B00",		-- 8, 11, 11, 8
        5949 => x"090B0B0B",		-- 9, 11, 11, 11
        5950 => x"0B0B0B09",		-- 11, 11, 11, 9
        5951 => x"000A0000",		-- 8, 10, 8, 8
        5952 => x"000B0B0A",		-- 8, 11, 11, 10
        5953 => x"0B0A090A",		-- 11, 10, 9, 10
        5954 => x"0B0B0B0B",		-- 11, 11, 11, 11
        5955 => x"000A0000",		-- 8, 10, 8, 8
        5956 => x"000B0B0A",		-- 8, 11, 11, 10
        5957 => x"0A0A0B0A",		-- 10, 10, 11, 10
        5958 => x"0A090A0B",		-- 10, 9, 10, 11
        5959 => x"0A0A0000",		-- 10, 10, 8, 8
        5960 => x"00000B0B",		-- 8, 8, 11, 11
        5961 => x"0A0A0A0A",		-- 10, 10, 10, 10
        5962 => x"0A0B0A0B",		-- 10, 11, 10, 11
        5963 => x"0A0A0000",		-- 10, 10, 8, 8
        5964 => x"00000B0B",		-- 8, 8, 11, 11
        5965 => x"0B0A0A0B",		-- 11, 10, 10, 11
        5966 => x"0A0A0A0A",		-- 10, 10, 10, 10
        5967 => x"0A0B0000",		-- 10, 11, 8, 8
        5968 => x"00000B0B",		-- 8, 8, 11, 11
        5969 => x"0B090A0B",		-- 11, 9, 10, 11
        5970 => x"0B0A0A09",		-- 11, 10, 10, 9
        5971 => x"0B0B0000",		-- 11, 11, 8, 8
        5972 => x"0000000B",		-- 8, 8, 8, 11
        5973 => x"09090909",		-- 9, 9, 9, 9
        5974 => x"0A0A0909",		-- 10, 10, 9, 9
        5975 => x"090A0000",		-- 9, 10, 8, 8
        5976 => x"0000000B",		-- 8, 8, 8, 11
        5977 => x"09090909",		-- 9, 9, 9, 9
        5978 => x"09090909",		-- 9, 9, 9, 9
        5979 => x"090A0000",		-- 9, 10, 8, 8
        5980 => x"00000009",		-- 8, 8, 8, 9
        5981 => x"09090B0B",		-- 9, 9, 11, 11
        5982 => x"0B0B0909",		-- 11, 11, 9, 9
        5983 => x"0B000000",		-- 11, 8, 8, 8
        5984 => x"0000000B",		-- 8, 8, 8, 11
        5985 => x"0B0B0B09",		-- 11, 11, 11, 9
        5986 => x"090B0B0B",		-- 9, 11, 11, 11
        5987 => x"09000000",		-- 9, 8, 8, 8
        5988 => x"00000009",		-- 8, 8, 8, 9
        5989 => x"09090B0B",		-- 9, 9, 11, 11
        5990 => x"0B0B0909",		-- 11, 11, 9, 9
        5991 => x"09000000",		-- 9, 8, 8, 8
        5992 => x"00000009",		-- 8, 8, 8, 9
        5993 => x"09090909",		-- 9, 9, 9, 9
        5994 => x"0909090B",		-- 9, 9, 9, 11
        5995 => x"00000000",		-- 8, 8, 8, 8
        5996 => x"00000000",		-- 8, 8, 8, 8
        5997 => x"0B0B0B00",		-- 11, 11, 11, 8
        5998 => x"000B0B0B",		-- 8, 11, 11, 11
        5999 => x"00000000",		-- 8, 8, 8, 8
        6000 => x"00000000",		-- 8, 8, 8, 8
        6001 => x"0B0B0B00",		-- 11, 11, 11, 8
        6002 => x"000B0B0B",		-- 8, 11, 11, 11
        6003 => x"00000000",		-- 8, 8, 8, 8

                --  sprite 13
        6004 => x"000A0A00",		-- 8, 10, 10, 8
        6005 => x"00000909",		-- 8, 8, 9, 9
        6006 => x"09090000",		-- 9, 9, 8, 8
        6007 => x"000A0A00",		-- 8, 10, 10, 8
        6008 => x"000A0A0A",		-- 8, 10, 10, 10
        6009 => x"00090B0B",		-- 8, 9, 11, 11
        6010 => x"0B0B0900",		-- 11, 11, 9, 8
        6011 => x"0A0A0A00",		-- 10, 10, 10, 8
        6012 => x"000B0B00",		-- 8, 11, 11, 8
        6013 => x"090B0B0B",		-- 9, 11, 11, 11
        6014 => x"0B0B0B09",		-- 11, 11, 11, 9
        6015 => x"000B0B00",		-- 8, 11, 11, 8
        6016 => x"000B0B0A",		-- 8, 11, 11, 10
        6017 => x"0B0A090A",		-- 11, 10, 9, 10
        6018 => x"0A090A0B",		-- 10, 9, 10, 11
        6019 => x"0A0B0B00",		-- 10, 11, 11, 8
        6020 => x"000B0B0A",		-- 8, 11, 11, 10
        6021 => x"0A0A0B0A",		-- 10, 10, 11, 10
        6022 => x"0A0B0A0A",		-- 10, 11, 10, 10
        6023 => x"0A0B0B00",		-- 10, 11, 11, 8
        6024 => x"00000B0B",		-- 8, 8, 11, 11
        6025 => x"0A0A0A0A",		-- 10, 10, 10, 10
        6026 => x"0A0A0A0A",		-- 10, 10, 10, 10
        6027 => x"0B0B0000",		-- 11, 11, 8, 8
        6028 => x"00000B0B",		-- 8, 8, 11, 11
        6029 => x"0B0A0A0B",		-- 11, 10, 10, 11
        6030 => x"0B0A0A0B",		-- 11, 10, 10, 11
        6031 => x"0B0B0000",		-- 11, 11, 8, 8
        6032 => x"00000B0B",		-- 8, 8, 11, 11
        6033 => x"0B090A0B",		-- 11, 9, 10, 11
        6034 => x"0B0A090B",		-- 11, 10, 9, 11
        6035 => x"0B0B0000",		-- 11, 11, 8, 8
        6036 => x"0000000B",		-- 8, 8, 8, 11
        6037 => x"09090909",		-- 9, 9, 9, 9
        6038 => x"09090909",		-- 9, 9, 9, 9
        6039 => x"0B000000",		-- 11, 8, 8, 8
        6040 => x"0000000B",		-- 8, 8, 8, 11
        6041 => x"09090909",		-- 9, 9, 9, 9
        6042 => x"09090909",		-- 9, 9, 9, 9
        6043 => x"0B000000",		-- 11, 8, 8, 8
        6044 => x"00000009",		-- 8, 8, 8, 9
        6045 => x"09090B0B",		-- 9, 9, 11, 11
        6046 => x"0B0B0909",		-- 11, 11, 9, 9
        6047 => x"09000000",		-- 9, 8, 8, 8
        6048 => x"0000000B",		-- 8, 8, 8, 11
        6049 => x"0B0B0B09",		-- 11, 11, 11, 9
        6050 => x"090B0B0B",		-- 9, 11, 11, 11
        6051 => x"0B000000",		-- 11, 8, 8, 8
        6052 => x"00000009",		-- 8, 8, 8, 9
        6053 => x"09090B0B",		-- 9, 9, 11, 11
        6054 => x"0B0B0909",		-- 11, 11, 9, 9
        6055 => x"09000000",		-- 9, 8, 8, 8
        6056 => x"00000009",		-- 8, 8, 8, 9
        6057 => x"09090909",		-- 9, 9, 9, 9
        6058 => x"09090909",		-- 9, 9, 9, 9
        6059 => x"09000000",		-- 9, 8, 8, 8
        6060 => x"00000000",		-- 8, 8, 8, 8
        6061 => x"0B0B0B00",		-- 11, 11, 11, 8
        6062 => x"000B0B0B",		-- 8, 11, 11, 11
        6063 => x"00000000",		-- 8, 8, 8, 8
        6064 => x"00000000",		-- 8, 8, 8, 8
        6065 => x"0B0B0B00",		-- 11, 11, 11, 8
        6066 => x"000B0B0B",		-- 8, 11, 11, 11
        6067 => x"00000000",		-- 8, 8, 8, 8

                --  sprite 14
        6068 => x"00000000",		-- 8, 8, 8, 8
        6069 => x"00000000",		-- 8, 8, 8, 8
        6070 => x"00000000",		-- 8, 8, 8, 8
        6071 => x"00000000",		-- 8, 8, 8, 8
        6072 => x"00000000",		-- 8, 8, 8, 8
        6073 => x"00000000",		-- 8, 8, 8, 8
        6074 => x"00000000",		-- 8, 8, 8, 8
        6075 => x"00000000",		-- 8, 8, 8, 8
        6076 => x"00000000",		-- 8, 8, 8, 8
        6077 => x"00000000",		-- 8, 8, 8, 8
        6078 => x"00000000",		-- 8, 8, 8, 8
        6079 => x"00000000",		-- 8, 8, 8, 8
        6080 => x"00000000",		-- 8, 8, 8, 8
        6081 => x"00000000",		-- 8, 8, 8, 8
        6082 => x"00000000",		-- 8, 8, 8, 8
        6083 => x"00000000",		-- 8, 8, 8, 8
        6084 => x"00000000",		-- 8, 8, 8, 8
        6085 => x"00000000",		-- 8, 8, 8, 8
        6086 => x"00000000",		-- 8, 8, 8, 8
        6087 => x"00000000",		-- 8, 8, 8, 8
        6088 => x"00000009",		-- 8, 8, 8, 9
        6089 => x"09000000",		-- 9, 8, 8, 8
        6090 => x"00000000",		-- 8, 8, 8, 8
        6091 => x"00000000",		-- 8, 8, 8, 8
        6092 => x"00000000",		-- 8, 8, 8, 8
        6093 => x"09000000",		-- 9, 8, 8, 8
        6094 => x"00000000",		-- 8, 8, 8, 8
        6095 => x"00000000",		-- 8, 8, 8, 8
        6096 => x"090A090A",		-- 9, 10, 9, 10
        6097 => x"090B0B0B",		-- 9, 11, 11, 11
        6098 => x"0B0B0B0B",		-- 11, 11, 11, 11
        6099 => x"0B0B0B00",		-- 11, 11, 11, 8
        6100 => x"090A090A",		-- 9, 10, 9, 10
        6101 => x"090B0B0B",		-- 9, 11, 11, 11
        6102 => x"0B0B0B0B",		-- 11, 11, 11, 11
        6103 => x"0B0B0B0B",		-- 11, 11, 11, 11
        6104 => x"090A090A",		-- 9, 10, 9, 10
        6105 => x"090B0B0B",		-- 9, 11, 11, 11
        6106 => x"0B0B0B0B",		-- 11, 11, 11, 11
        6107 => x"0B0B0B00",		-- 11, 11, 11, 8
        6108 => x"00000000",		-- 8, 8, 8, 8
        6109 => x"09000000",		-- 9, 8, 8, 8
        6110 => x"00000000",		-- 8, 8, 8, 8
        6111 => x"00000000",		-- 8, 8, 8, 8
        6112 => x"00000009",		-- 8, 8, 8, 9
        6113 => x"09000000",		-- 9, 8, 8, 8
        6114 => x"00000000",		-- 8, 8, 8, 8
        6115 => x"00000000",		-- 8, 8, 8, 8
        6116 => x"00000000",		-- 8, 8, 8, 8
        6117 => x"00000000",		-- 8, 8, 8, 8
        6118 => x"00000000",		-- 8, 8, 8, 8
        6119 => x"00000000",		-- 8, 8, 8, 8
        6120 => x"00000000",		-- 8, 8, 8, 8
        6121 => x"00000000",		-- 8, 8, 8, 8
        6122 => x"00000000",		-- 8, 8, 8, 8
        6123 => x"00000000",		-- 8, 8, 8, 8
        6124 => x"00000000",		-- 8, 8, 8, 8
        6125 => x"00000000",		-- 8, 8, 8, 8
        6126 => x"00000000",		-- 8, 8, 8, 8
        6127 => x"00000000",		-- 8, 8, 8, 8
        6128 => x"00000000",		-- 8, 8, 8, 8
        6129 => x"00000000",		-- 8, 8, 8, 8
        6130 => x"00000000",		-- 8, 8, 8, 8
        6131 => x"00000000",		-- 8, 8, 8, 8

                --  sprite 15
        6132 => x"00000000",		-- 8, 8, 8, 8
        6133 => x"00000000",		-- 8, 8, 8, 8
        6134 => x"00000000",		-- 8, 8, 8, 8
        6135 => x"00000000",		-- 8, 8, 8, 8
        6136 => x"00000000",		-- 8, 8, 8, 8
        6137 => x"00000000",		-- 8, 8, 8, 8
        6138 => x"00000000",		-- 8, 8, 8, 8
        6139 => x"00000000",		-- 8, 8, 8, 8
        6140 => x"00000000",		-- 8, 8, 8, 8
        6141 => x"00000000",		-- 8, 8, 8, 8
        6142 => x"00000000",		-- 8, 8, 8, 8
        6143 => x"00000000",		-- 8, 8, 8, 8
        6144 => x"00000000",		-- 8, 8, 8, 8
        6145 => x"00000000",		-- 8, 8, 8, 8
        6146 => x"00000000",		-- 8, 8, 8, 8
        6147 => x"00000000",		-- 8, 8, 8, 8
        6148 => x"00000000",		-- 8, 8, 8, 8
        6149 => x"00000000",		-- 8, 8, 8, 8
        6150 => x"00000000",		-- 8, 8, 8, 8
        6151 => x"00000000",		-- 8, 8, 8, 8
        6152 => x"0B000B00",		-- 11, 8, 11, 8
        6153 => x"0B000000",		-- 11, 8, 8, 8
        6154 => x"00000000",		-- 8, 8, 8, 8
        6155 => x"00000000",		-- 8, 8, 8, 8
        6156 => x"000B000B",		-- 8, 11, 8, 11
        6157 => x"000B0000",		-- 8, 11, 8, 8
        6158 => x"00000000",		-- 8, 8, 8, 8
        6159 => x"0A0A0000",		-- 10, 10, 8, 8
        6160 => x"09090909",		-- 9, 9, 9, 9
        6161 => x"09090909",		-- 9, 9, 9, 9
        6162 => x"09090909",		-- 9, 9, 9, 9
        6163 => x"090A0A0A",		-- 9, 10, 10, 10
        6164 => x"000B000B",		-- 8, 11, 8, 11
        6165 => x"000B0000",		-- 8, 11, 8, 8
        6166 => x"00000000",		-- 8, 8, 8, 8
        6167 => x"0A0A0000",		-- 10, 10, 8, 8
        6168 => x"0B000B00",		-- 11, 8, 11, 8
        6169 => x"0B000000",		-- 11, 8, 8, 8
        6170 => x"00000000",		-- 8, 8, 8, 8
        6171 => x"00000000",		-- 8, 8, 8, 8
        6172 => x"00000000",		-- 8, 8, 8, 8
        6173 => x"00000000",		-- 8, 8, 8, 8
        6174 => x"00000000",		-- 8, 8, 8, 8
        6175 => x"00000000",		-- 8, 8, 8, 8
        6176 => x"00000000",		-- 8, 8, 8, 8
        6177 => x"00000000",		-- 8, 8, 8, 8
        6178 => x"00000000",		-- 8, 8, 8, 8
        6179 => x"00000000",		-- 8, 8, 8, 8
        6180 => x"00000000",		-- 8, 8, 8, 8
        6181 => x"00000000",		-- 8, 8, 8, 8
        6182 => x"00000000",		-- 8, 8, 8, 8
        6183 => x"00000000",		-- 8, 8, 8, 8
        6184 => x"00000000",		-- 8, 8, 8, 8
        6185 => x"00000000",		-- 8, 8, 8, 8
        6186 => x"00000000",		-- 8, 8, 8, 8
        6187 => x"00000000",		-- 8, 8, 8, 8
        6188 => x"00000000",		-- 8, 8, 8, 8
        6189 => x"00000000",		-- 8, 8, 8, 8
        6190 => x"00000000",		-- 8, 8, 8, 8
        6191 => x"00000000",		-- 8, 8, 8, 8
        6192 => x"00000000",		-- 8, 8, 8, 8
        6193 => x"00000000",		-- 8, 8, 8, 8
        6194 => x"00000000",		-- 8, 8, 8, 8
        6195 => x"00000000",		-- 8, 8, 8, 8

                --  sprite 16
        6196 => x"00000000",		-- 8, 8, 8, 8
        6197 => x"00000000",		-- 8, 8, 8, 8
        6198 => x"12121212",		-- 18, 18, 18, 18
        6199 => x"12121212",		-- 18, 18, 18, 18
        6200 => x"00000000",		-- 8, 8, 8, 8
        6201 => x"00000000",		-- 8, 8, 8, 8
        6202 => x"12121212",		-- 18, 18, 18, 18
        6203 => x"12121212",		-- 18, 18, 18, 18
        6204 => x"00000000",		-- 8, 8, 8, 8
        6205 => x"00000000",		-- 8, 8, 8, 8
        6206 => x"12121212",		-- 18, 18, 18, 18
        6207 => x"12121212",		-- 18, 18, 18, 18
        6208 => x"00000000",		-- 8, 8, 8, 8
        6209 => x"00000000",		-- 8, 8, 8, 8
        6210 => x"12121212",		-- 18, 18, 18, 18
        6211 => x"12121212",		-- 18, 18, 18, 18
        6212 => x"0A0B0000",		-- 10, 11, 8, 8
        6213 => x"00000000",		-- 8, 8, 8, 8
        6214 => x"12121212",		-- 18, 18, 18, 18
        6215 => x"12121212",		-- 18, 18, 18, 18
        6216 => x"0A0B0000",		-- 10, 11, 8, 8
        6217 => x"00000000",		-- 8, 8, 8, 8
        6218 => x"12121212",		-- 18, 18, 18, 18
        6219 => x"12121212",		-- 18, 18, 18, 18
        6220 => x"0A090B00",		-- 10, 9, 11, 8
        6221 => x"00000000",		-- 8, 8, 8, 8
        6222 => x"12121212",		-- 18, 18, 18, 18
        6223 => x"12121212",		-- 18, 18, 18, 18
        6224 => x"0909090B",		-- 9, 9, 9, 11
        6225 => x"00000000",		-- 8, 8, 8, 8
        6226 => x"12121212",		-- 18, 18, 18, 18
        6227 => x"12121212",		-- 18, 18, 18, 18
        6228 => x"00090A0A",		-- 8, 9, 10, 10
        6229 => x"0B000000",		-- 11, 8, 8, 8
        6230 => x"12121212",		-- 18, 18, 18, 18
        6231 => x"12121212",		-- 18, 18, 18, 18
        6232 => x"000A0A0A",		-- 8, 10, 10, 10
        6233 => x"0A0B0000",		-- 10, 11, 8, 8
        6234 => x"12121212",		-- 18, 18, 18, 18
        6235 => x"12121212",		-- 18, 18, 18, 18
        6236 => x"00000A0A",		-- 8, 8, 10, 10
        6237 => x"0A0A0B0B",		-- 10, 10, 11, 11
        6238 => x"12121212",		-- 18, 18, 18, 18
        6239 => x"12121212",		-- 18, 18, 18, 18
        6240 => x"00000000",		-- 8, 8, 8, 8
        6241 => x"0A0A0A0A",		-- 10, 10, 10, 10
        6242 => x"12121212",		-- 18, 18, 18, 18
        6243 => x"12121212",		-- 18, 18, 18, 18
        6244 => x"00000000",		-- 8, 8, 8, 8
        6245 => x"00000000",		-- 8, 8, 8, 8
        6246 => x"12121212",		-- 18, 18, 18, 18
        6247 => x"12121212",		-- 18, 18, 18, 18
        6248 => x"00000000",		-- 8, 8, 8, 8
        6249 => x"00000000",		-- 8, 8, 8, 8
        6250 => x"12121212",		-- 18, 18, 18, 18
        6251 => x"12121212",		-- 18, 18, 18, 18
        6252 => x"00000000",		-- 8, 8, 8, 8
        6253 => x"00000000",		-- 8, 8, 8, 8
        6254 => x"12121212",		-- 18, 18, 18, 18
        6255 => x"12121212",		-- 18, 18, 18, 18
        6256 => x"00000000",		-- 8, 8, 8, 8
        6257 => x"00000000",		-- 8, 8, 8, 8
        6258 => x"12121212",		-- 18, 18, 18, 18
        6259 => x"12121212",		-- 18, 18, 18, 18

                --  sprite 17
        6260 => x"00000000",		-- 8, 8, 8, 8
        6261 => x"00000000",		-- 8, 8, 8, 8
        6262 => x"12121212",		-- 18, 18, 18, 18
        6263 => x"12121212",		-- 18, 18, 18, 18
        6264 => x"00000000",		-- 8, 8, 8, 8
        6265 => x"00000000",		-- 8, 8, 8, 8
        6266 => x"12121212",		-- 18, 18, 18, 18
        6267 => x"12121212",		-- 18, 18, 18, 18
        6268 => x"00000000",		-- 8, 8, 8, 8
        6269 => x"00000000",		-- 8, 8, 8, 8
        6270 => x"12121212",		-- 18, 18, 18, 18
        6271 => x"12121212",		-- 18, 18, 18, 18
        6272 => x"00000000",		-- 8, 8, 8, 8
        6273 => x"00000000",		-- 8, 8, 8, 8
        6274 => x"12121212",		-- 18, 18, 18, 18
        6275 => x"12121212",		-- 18, 18, 18, 18
        6276 => x"00000000",		-- 8, 8, 8, 8
        6277 => x"00000000",		-- 8, 8, 8, 8
        6278 => x"12121212",		-- 18, 18, 18, 18
        6279 => x"12121212",		-- 18, 18, 18, 18
        6280 => x"00000000",		-- 8, 8, 8, 8
        6281 => x"00000000",		-- 8, 8, 8, 8
        6282 => x"12121212",		-- 18, 18, 18, 18
        6283 => x"12121212",		-- 18, 18, 18, 18
        6284 => x"0B000000",		-- 11, 8, 8, 8
        6285 => x"0000000B",		-- 8, 8, 8, 11
        6286 => x"12121212",		-- 18, 18, 18, 18
        6287 => x"12121212",		-- 18, 18, 18, 18
        6288 => x"0A0B0000",		-- 10, 11, 8, 8
        6289 => x"00000B0A",		-- 8, 8, 11, 10
        6290 => x"12121212",		-- 18, 18, 18, 18
        6291 => x"12121212",		-- 18, 18, 18, 18
        6292 => x"09090B0B",		-- 9, 9, 11, 11
        6293 => x"0B0B0A0A",		-- 11, 11, 10, 10
        6294 => x"12121212",		-- 18, 18, 18, 18
        6295 => x"12121212",		-- 18, 18, 18, 18
        6296 => x"0009090A",		-- 8, 9, 9, 10
        6297 => x"0A0A0A00",		-- 10, 10, 10, 8
        6298 => x"12121212",		-- 18, 18, 18, 18
        6299 => x"12121212",		-- 18, 18, 18, 18
        6300 => x"00000A0A",		-- 8, 8, 10, 10
        6301 => x"0A0A0000",		-- 10, 10, 8, 8
        6302 => x"12121212",		-- 18, 18, 18, 18
        6303 => x"12121212",		-- 18, 18, 18, 18
        6304 => x"00000000",		-- 8, 8, 8, 8
        6305 => x"00000000",		-- 8, 8, 8, 8
        6306 => x"12121212",		-- 18, 18, 18, 18
        6307 => x"12121212",		-- 18, 18, 18, 18
        6308 => x"00000000",		-- 8, 8, 8, 8
        6309 => x"00000000",		-- 8, 8, 8, 8
        6310 => x"12121212",		-- 18, 18, 18, 18
        6311 => x"12121212",		-- 18, 18, 18, 18
        6312 => x"00000000",		-- 8, 8, 8, 8
        6313 => x"00000000",		-- 8, 8, 8, 8
        6314 => x"12121212",		-- 18, 18, 18, 18
        6315 => x"12121212",		-- 18, 18, 18, 18
        6316 => x"00000000",		-- 8, 8, 8, 8
        6317 => x"00000000",		-- 8, 8, 8, 8
        6318 => x"12121212",		-- 18, 18, 18, 18
        6319 => x"12121212",		-- 18, 18, 18, 18
        6320 => x"00000000",		-- 8, 8, 8, 8
        6321 => x"00000000",		-- 8, 8, 8, 8
        6322 => x"12121212",		-- 18, 18, 18, 18
        6323 => x"12121212",		-- 18, 18, 18, 18

                --  sprite 18
        6324 => x"00000000",		-- 8, 8, 8, 8
        6325 => x"00090909",		-- 8, 9, 9, 9
        6326 => x"09090900",		-- 9, 9, 9, 8
        6327 => x"00000000",		-- 8, 8, 8, 8
        6328 => x"00000009",		-- 8, 8, 8, 9
        6329 => x"09090909",		-- 9, 9, 9, 9
        6330 => x"09090909",		-- 9, 9, 9, 9
        6331 => x"09000000",		-- 9, 8, 8, 8
        6332 => x"00000909",		-- 8, 8, 9, 9
        6333 => x"09090909",		-- 9, 9, 9, 9
        6334 => x"09090909",		-- 9, 9, 9, 9
        6335 => x"09090000",		-- 9, 9, 8, 8
        6336 => x"00090909",		-- 8, 9, 9, 9
        6337 => x"00000000",		-- 8, 8, 8, 8
        6338 => x"00000000",		-- 8, 8, 8, 8
        6339 => x"09090900",		-- 9, 9, 9, 8
        6340 => x"00090000",		-- 8, 9, 8, 8
        6341 => x"00000000",		-- 8, 8, 8, 8
        6342 => x"00000000",		-- 8, 8, 8, 8
        6343 => x"00000900",		-- 8, 8, 9, 8
        6344 => x"09000000",		-- 9, 8, 8, 8
        6345 => x"000A0A0A",		-- 8, 10, 10, 10
        6346 => x"0A0A0A00",		-- 10, 10, 10, 8
        6347 => x"00000009",		-- 8, 8, 8, 9
        6348 => x"0000000A",		-- 8, 8, 8, 10
        6349 => x"0A0A0A0A",		-- 10, 10, 10, 10
        6350 => x"0A0A0A0A",		-- 10, 10, 10, 10
        6351 => x"0A000000",		-- 10, 8, 8, 8
        6352 => x"00000A0A",		-- 8, 8, 10, 10
        6353 => x"0A0A0000",		-- 10, 10, 8, 8
        6354 => x"00000A0A",		-- 8, 8, 10, 10
        6355 => x"0A0A0000",		-- 10, 10, 8, 8
        6356 => x"000A0A00",		-- 8, 10, 10, 8
        6357 => x"00000000",		-- 8, 8, 8, 8
        6358 => x"00000000",		-- 8, 8, 8, 8
        6359 => x"000A0A00",		-- 8, 10, 10, 8
        6360 => x"000A0000",		-- 8, 10, 8, 8
        6361 => x"00000909",		-- 8, 8, 9, 9
        6362 => x"09090000",		-- 9, 9, 8, 8
        6363 => x"00000A00",		-- 8, 8, 10, 8
        6364 => x"00000000",		-- 8, 8, 8, 8
        6365 => x"09090909",		-- 9, 9, 9, 9
        6366 => x"09090909",		-- 9, 9, 9, 9
        6367 => x"00000000",		-- 8, 8, 8, 8
        6368 => x"00000009",		-- 8, 8, 8, 9
        6369 => x"09000000",		-- 9, 8, 8, 8
        6370 => x"00000009",		-- 8, 8, 8, 9
        6371 => x"09000000",		-- 9, 8, 8, 8
        6372 => x"00000900",		-- 8, 8, 9, 8
        6373 => x"0000000A",		-- 8, 8, 8, 10
        6374 => x"0A000000",		-- 10, 8, 8, 8
        6375 => x"00090000",		-- 8, 9, 8, 8
        6376 => x"00000000",		-- 8, 8, 8, 8
        6377 => x"000A0A0A",		-- 8, 10, 10, 10
        6378 => x"0A0A0A00",		-- 10, 10, 10, 8
        6379 => x"00000000",		-- 8, 8, 8, 8
        6380 => x"00000000",		-- 8, 8, 8, 8
        6381 => x"0A0A0000",		-- 10, 10, 8, 8
        6382 => x"00000A0A",		-- 8, 8, 10, 10
        6383 => x"00000000",		-- 8, 8, 8, 8
        6384 => x"0000000A",		-- 8, 8, 8, 10
        6385 => x"00000000",		-- 8, 8, 8, 8
        6386 => x"00000000",		-- 8, 8, 8, 8
        6387 => x"0A000000",		-- 10, 8, 8, 8

                --  sprite 19
        6388 => x"00000000",		-- 8, 8, 8, 8
        6389 => x"00000000",		-- 8, 8, 8, 8
        6390 => x"00000900",		-- 8, 8, 9, 8
        6391 => x"00000000",		-- 8, 8, 8, 8
        6392 => x"00000000",		-- 8, 8, 8, 8
        6393 => x"00000A0A",		-- 8, 8, 10, 10
        6394 => x"00000009",		-- 8, 8, 8, 9
        6395 => x"09000000",		-- 9, 8, 8, 8
        6396 => x"00000009",		-- 8, 8, 8, 9
        6397 => x"0000000A",		-- 8, 8, 8, 10
        6398 => x"0A000000",		-- 10, 8, 8, 8
        6399 => x"09090000",		-- 9, 9, 8, 8
        6400 => x"0A000000",		-- 10, 8, 8, 8
        6401 => x"09000000",		-- 9, 8, 8, 8
        6402 => x"0A0A0000",		-- 10, 10, 8, 8
        6403 => x"09090900",		-- 9, 9, 9, 8
        6404 => x"000A0000",		-- 8, 10, 8, 8
        6405 => x"09090000",		-- 9, 9, 8, 8
        6406 => x"0A0A0000",		-- 10, 10, 8, 8
        6407 => x"00090900",		-- 8, 9, 9, 8
        6408 => x"000A0A00",		-- 8, 10, 10, 8
        6409 => x"00090000",		-- 8, 9, 8, 8
        6410 => x"0A0A0A00",		-- 10, 10, 10, 8
        6411 => x"00090909",		-- 8, 9, 9, 9
        6412 => x"00000A00",		-- 8, 8, 10, 8
        6413 => x"00090900",		-- 8, 9, 9, 8
        6414 => x"000A0A00",		-- 8, 10, 10, 8
        6415 => x"00090909",		-- 8, 9, 9, 9
        6416 => x"00000A0A",		-- 8, 8, 10, 10
        6417 => x"00090900",		-- 8, 9, 9, 8
        6418 => x"000A0A00",		-- 8, 10, 10, 8
        6419 => x"00090909",		-- 8, 9, 9, 9
        6420 => x"00000A0A",		-- 8, 8, 10, 10
        6421 => x"00090900",		-- 8, 9, 9, 8
        6422 => x"000A0A00",		-- 8, 10, 10, 8
        6423 => x"00090909",		-- 8, 9, 9, 9
        6424 => x"00000A00",		-- 8, 8, 10, 8
        6425 => x"00090900",		-- 8, 9, 9, 8
        6426 => x"000A0A00",		-- 8, 10, 10, 8
        6427 => x"00090909",		-- 8, 9, 9, 9
        6428 => x"000A0A00",		-- 8, 10, 10, 8
        6429 => x"00090000",		-- 8, 9, 8, 8
        6430 => x"0A0A0A00",		-- 10, 10, 10, 8
        6431 => x"00090909",		-- 8, 9, 9, 9
        6432 => x"000A0000",		-- 8, 10, 8, 8
        6433 => x"09090000",		-- 9, 9, 8, 8
        6434 => x"0A0A0000",		-- 10, 10, 8, 8
        6435 => x"00090900",		-- 8, 9, 9, 8
        6436 => x"0A000000",		-- 10, 8, 8, 8
        6437 => x"09000000",		-- 9, 8, 8, 8
        6438 => x"0A0A0000",		-- 10, 10, 8, 8
        6439 => x"09090900",		-- 9, 9, 9, 8
        6440 => x"00000009",		-- 8, 8, 8, 9
        6441 => x"0000000A",		-- 8, 8, 8, 10
        6442 => x"0A000000",		-- 10, 8, 8, 8
        6443 => x"09090000",		-- 9, 9, 8, 8
        6444 => x"00000000",		-- 8, 8, 8, 8
        6445 => x"00000A0A",		-- 8, 8, 10, 10
        6446 => x"00000009",		-- 8, 8, 8, 9
        6447 => x"09000000",		-- 9, 8, 8, 8
        6448 => x"00000000",		-- 8, 8, 8, 8
        6449 => x"00000000",		-- 8, 8, 8, 8
        6450 => x"00000900",		-- 8, 8, 9, 8
        6451 => x"00000000",		-- 8, 8, 8, 8

                --  sprite 20
        6452 => x"00000000",		-- 8, 8, 8, 8
        6453 => x"00000000",		-- 8, 8, 8, 8
        6454 => x"12121212",		-- 18, 18, 18, 18
        6455 => x"12121212",		-- 18, 18, 18, 18
        6456 => x"00000000",		-- 8, 8, 8, 8
        6457 => x"00000000",		-- 8, 8, 8, 8
        6458 => x"12121212",		-- 18, 18, 18, 18
        6459 => x"12121212",		-- 18, 18, 18, 18
        6460 => x"00000000",		-- 8, 8, 8, 8
        6461 => x"00000000",		-- 8, 8, 8, 8
        6462 => x"12121212",		-- 18, 18, 18, 18
        6463 => x"12121212",		-- 18, 18, 18, 18
        6464 => x"00000000",		-- 8, 8, 8, 8
        6465 => x"00000000",		-- 8, 8, 8, 8
        6466 => x"12121212",		-- 18, 18, 18, 18
        6467 => x"12121212",		-- 18, 18, 18, 18
        6468 => x"000F0000",		-- 8, 15, 8, 8
        6469 => x"000F0000",		-- 8, 15, 8, 8
        6470 => x"12121212",		-- 18, 18, 18, 18
        6471 => x"12121212",		-- 18, 18, 18, 18
        6472 => x"00000F00",		-- 8, 8, 15, 8
        6473 => x"0F0F000F",		-- 15, 15, 8, 15
        6474 => x"12121212",		-- 18, 18, 18, 18
        6475 => x"12121212",		-- 18, 18, 18, 18
        6476 => x"0F000F0F",		-- 15, 8, 15, 15
        6477 => x"0F0F0F00",		-- 15, 15, 15, 8
        6478 => x"12121212",		-- 18, 18, 18, 18
        6479 => x"12121212",		-- 18, 18, 18, 18
        6480 => x"000F0F0F",		-- 8, 15, 15, 15
        6481 => x"0F0F0000",		-- 15, 15, 8, 8
        6482 => x"12121212",		-- 18, 18, 18, 18
        6483 => x"12121212",		-- 18, 18, 18, 18
        6484 => x"00000F0F",		-- 8, 8, 15, 15
        6485 => x"0F000000",		-- 15, 8, 8, 8
        6486 => x"12121212",		-- 18, 18, 18, 18
        6487 => x"12121212",		-- 18, 18, 18, 18
        6488 => x"000F0F0F",		-- 8, 15, 15, 15
        6489 => x"0F0F0000",		-- 15, 15, 8, 8
        6490 => x"12121212",		-- 18, 18, 18, 18
        6491 => x"12121212",		-- 18, 18, 18, 18
        6492 => x"0F00000F",		-- 15, 8, 8, 15
        6493 => x"00000000",		-- 8, 8, 8, 8
        6494 => x"12121212",		-- 18, 18, 18, 18
        6495 => x"12121212",		-- 18, 18, 18, 18
        6496 => x"00000000",		-- 8, 8, 8, 8
        6497 => x"0F000000",		-- 15, 8, 8, 8
        6498 => x"12121212",		-- 18, 18, 18, 18
        6499 => x"12121212",		-- 18, 18, 18, 18
        6500 => x"00000000",		-- 8, 8, 8, 8
        6501 => x"00000000",		-- 8, 8, 8, 8
        6502 => x"12121212",		-- 18, 18, 18, 18
        6503 => x"12121212",		-- 18, 18, 18, 18
        6504 => x"00000000",		-- 8, 8, 8, 8
        6505 => x"00000000",		-- 8, 8, 8, 8
        6506 => x"12121212",		-- 18, 18, 18, 18
        6507 => x"12121212",		-- 18, 18, 18, 18
        6508 => x"00000000",		-- 8, 8, 8, 8
        6509 => x"00000000",		-- 8, 8, 8, 8
        6510 => x"12121212",		-- 18, 18, 18, 18
        6511 => x"12121212",		-- 18, 18, 18, 18
        6512 => x"00000000",		-- 8, 8, 8, 8
        6513 => x"00000000",		-- 8, 8, 8, 8
        6514 => x"12121212",		-- 18, 18, 18, 18
        6515 => x"12121212",		-- 18, 18, 18, 18

                --  sprite 21
        6516 => x"00000000",		-- 8, 8, 8, 8
        6517 => x"00090909",		-- 8, 9, 9, 9
        6518 => x"09090900",		-- 9, 9, 9, 8
        6519 => x"00000000",		-- 8, 8, 8, 8
        6520 => x"00000000",		-- 8, 8, 8, 8
        6521 => x"09090909",		-- 9, 9, 9, 9
        6522 => x"09090909",		-- 9, 9, 9, 9
        6523 => x"00000000",		-- 8, 8, 8, 8
        6524 => x"00000A00",		-- 8, 8, 10, 8
        6525 => x"09090909",		-- 9, 9, 9, 9
        6526 => x"09090909",		-- 9, 9, 9, 9
        6527 => x"000A0000",		-- 8, 10, 8, 8
        6528 => x"00000A09",		-- 8, 8, 10, 9
        6529 => x"09090909",		-- 9, 9, 9, 9
        6530 => x"09090909",		-- 9, 9, 9, 9
        6531 => x"090A0000",		-- 9, 10, 8, 8
        6532 => x"00000A0B",		-- 8, 8, 10, 11
        6533 => x"09090909",		-- 9, 9, 9, 9
        6534 => x"09090909",		-- 9, 9, 9, 9
        6535 => x"0B0A0000",		-- 11, 10, 8, 8
        6536 => x"00000A0A",		-- 8, 8, 10, 10
        6537 => x"0B0B0909",		-- 11, 11, 9, 9
        6538 => x"09090B0B",		-- 9, 9, 11, 11
        6539 => x"0A0A0000",		-- 10, 10, 8, 8
        6540 => x"0000000A",		-- 8, 8, 8, 10
        6541 => x"0B0B0B09",		-- 11, 11, 11, 9
        6542 => x"090B0B0B",		-- 9, 11, 11, 11
        6543 => x"0A000000",		-- 10, 8, 8, 8
        6544 => x"0000000B",		-- 8, 8, 8, 11
        6545 => x"090B0B0B",		-- 9, 11, 11, 11
        6546 => x"0B0B0B09",		-- 11, 11, 11, 9
        6547 => x"0B000000",		-- 11, 8, 8, 8
        6548 => x"00000B0B",		-- 8, 8, 11, 11
        6549 => x"09090909",		-- 9, 9, 9, 9
        6550 => x"0909090B",		-- 9, 9, 9, 11
        6551 => x"0B000000",		-- 11, 8, 8, 8
        6552 => x"00000B0B",		-- 8, 8, 11, 11
        6553 => x"09090909",		-- 9, 9, 9, 9
        6554 => x"0909090B",		-- 9, 9, 9, 11
        6555 => x"0B0A0000",		-- 11, 10, 8, 8
        6556 => x"0000000B",		-- 8, 8, 8, 11
        6557 => x"0B090909",		-- 11, 9, 9, 9
        6558 => x"0909090B",		-- 9, 9, 9, 11
        6559 => x"0B0A0000",		-- 11, 10, 8, 8
        6560 => x"00000009",		-- 8, 8, 8, 9
        6561 => x"090B0B0B",		-- 9, 11, 11, 11
        6562 => x"0B0B0B09",		-- 11, 11, 11, 9
        6563 => x"0A0A0000",		-- 10, 10, 8, 8
        6564 => x"00000009",		-- 8, 8, 8, 9
        6565 => x"09090909",		-- 9, 9, 9, 9
        6566 => x"09090909",		-- 9, 9, 9, 9
        6567 => x"09000000",		-- 9, 8, 8, 8
        6568 => x"0000000B",		-- 8, 8, 8, 11
        6569 => x"0B0B0909",		-- 11, 11, 9, 9
        6570 => x"0909090B",		-- 9, 9, 9, 11
        6571 => x"00000000",		-- 8, 8, 8, 8
        6572 => x"0000000B",		-- 8, 8, 8, 11
        6573 => x"0B0B0B00",		-- 11, 11, 11, 8
        6574 => x"000B0B00",		-- 8, 11, 11, 8
        6575 => x"00000000",		-- 8, 8, 8, 8
        6576 => x"00000000",		-- 8, 8, 8, 8
        6577 => x"0B0B0000",		-- 11, 11, 8, 8
        6578 => x"00000000",		-- 8, 8, 8, 8
        6579 => x"00000000",		-- 8, 8, 8, 8

                --  sprite 22
        6580 => x"00000000",		-- 8, 8, 8, 8
        6581 => x"00000000",		-- 8, 8, 8, 8
        6582 => x"00000000",		-- 8, 8, 8, 8
        6583 => x"00000000",		-- 8, 8, 8, 8
        6584 => x"00000000",		-- 8, 8, 8, 8
        6585 => x"00000009",		-- 8, 8, 8, 9
        6586 => x"09090900",		-- 9, 9, 9, 8
        6587 => x"00000000",		-- 8, 8, 8, 8
        6588 => x"00000000",		-- 8, 8, 8, 8
        6589 => x"0B0B0B0B",		-- 11, 11, 11, 11
        6590 => x"09090909",		-- 9, 9, 9, 9
        6591 => x"09000000",		-- 9, 8, 8, 8
        6592 => x"0000000B",		-- 8, 8, 8, 11
        6593 => x"0B0B0B0B",		-- 11, 11, 11, 11
        6594 => x"0B09090A",		-- 11, 9, 9, 10
        6595 => x"09090900",		-- 9, 9, 9, 8
        6596 => x"00000000",		-- 8, 8, 8, 8
        6597 => x"0B0B0B0B",		-- 11, 11, 11, 11
        6598 => x"0B0B0A0A",		-- 11, 11, 10, 10
        6599 => x"09090909",		-- 9, 9, 9, 9
        6600 => x"00000000",		-- 8, 8, 8, 8
        6601 => x"0A090A0A",		-- 10, 9, 10, 10
        6602 => x"0B0A0A0A",		-- 11, 10, 10, 10
        6603 => x"09090009",		-- 9, 9, 8, 9
        6604 => x"00000A0A",		-- 8, 8, 10, 10
        6605 => x"0A0B0A0A",		-- 10, 11, 10, 10
        6606 => x"0B0A0A0B",		-- 11, 10, 10, 11
        6607 => x"0B090000",		-- 11, 9, 8, 8
        6608 => x"00000B00",		-- 8, 8, 11, 8
        6609 => x"0A0A0A0A",		-- 10, 10, 10, 10
        6610 => x"0A0A0B0B",		-- 10, 10, 11, 11
        6611 => x"0B000000",		-- 11, 8, 8, 8
        6612 => x"00000B00",		-- 8, 8, 11, 8
        6613 => x"0A0A0A0A",		-- 10, 10, 10, 10
        6614 => x"09090909",		-- 9, 9, 9, 9
        6615 => x"00000000",		-- 8, 8, 8, 8
        6616 => x"00000B0A",		-- 8, 8, 11, 10
        6617 => x"0B0B0A0A",		-- 11, 11, 10, 10
        6618 => x"0A09090B",		-- 10, 9, 9, 11
        6619 => x"0B090000",		-- 11, 9, 8, 8
        6620 => x"00000B0A",		-- 8, 8, 11, 10
        6621 => x"0B090A0A",		-- 11, 9, 10, 10
        6622 => x"0A0B0B0B",		-- 10, 11, 11, 11
        6623 => x"0B0B0000",		-- 11, 11, 8, 8
        6624 => x"00000B00",		-- 8, 8, 11, 8
        6625 => x"0B09090A",		-- 11, 9, 9, 10
        6626 => x"0A0B0B0B",		-- 10, 11, 11, 11
        6627 => x"0B0B0900",		-- 11, 11, 9, 8
        6628 => x"00000B00",		-- 8, 8, 11, 8
        6629 => x"000B0909",		-- 8, 11, 9, 9
        6630 => x"090B0B0B",		-- 9, 11, 11, 11
        6631 => x"0B090900",		-- 11, 9, 9, 8
        6632 => x"00000B00",		-- 8, 8, 11, 8
        6633 => x"090B0B0B",		-- 9, 11, 11, 11
        6634 => x"0B090909",		-- 11, 9, 9, 9
        6635 => x"09090B0B",		-- 9, 9, 11, 11
        6636 => x"0000000B",		-- 8, 8, 8, 11
        6637 => x"0B090909",		-- 11, 9, 9, 9
        6638 => x"09090909",		-- 9, 9, 9, 9
        6639 => x"090B0B0B",		-- 9, 11, 11, 11
        6640 => x"00000000",		-- 8, 8, 8, 8
        6641 => x"0B0B0B00",		-- 11, 11, 11, 8
        6642 => x"00000000",		-- 8, 8, 8, 8
        6643 => x"0B0B0B00",		-- 11, 11, 11, 8

                --  sprite 23
        6644 => x"00000000",		-- 8, 8, 8, 8
        6645 => x"00000009",		-- 8, 8, 8, 9
        6646 => x"09090900",		-- 9, 9, 9, 8
        6647 => x"00000000",		-- 8, 8, 8, 8
        6648 => x"00000000",		-- 8, 8, 8, 8
        6649 => x"0B0B0B0B",		-- 11, 11, 11, 11
        6650 => x"09090909",		-- 9, 9, 9, 9
        6651 => x"09000000",		-- 9, 8, 8, 8
        6652 => x"0000000B",		-- 8, 8, 8, 11
        6653 => x"0B0B0B0B",		-- 11, 11, 11, 11
        6654 => x"0B09090A",		-- 11, 9, 9, 10
        6655 => x"09090900",		-- 9, 9, 9, 8
        6656 => x"00000000",		-- 8, 8, 8, 8
        6657 => x"0B0B0B0B",		-- 11, 11, 11, 11
        6658 => x"0B0B0A0A",		-- 11, 11, 10, 10
        6659 => x"09090909",		-- 9, 9, 9, 9
        6660 => x"000B0000",		-- 8, 11, 8, 8
        6661 => x"0A090A0A",		-- 10, 9, 10, 10
        6662 => x"0B0A0A0A",		-- 11, 10, 10, 10
        6663 => x"09090009",		-- 9, 9, 8, 9
        6664 => x"000B0A0A",		-- 8, 11, 10, 10
        6665 => x"0A0B0A0A",		-- 10, 11, 10, 10
        6666 => x"0B0A0A0B",		-- 11, 10, 10, 11
        6667 => x"0B090000",		-- 11, 9, 8, 8
        6668 => x"000B0000",		-- 8, 11, 8, 8
        6669 => x"0A0A0A0A",		-- 10, 10, 10, 10
        6670 => x"0A0A0B0B",		-- 10, 10, 11, 11
        6671 => x"0B000000",		-- 11, 8, 8, 8
        6672 => x"000B0000",		-- 8, 11, 8, 8
        6673 => x"0A0A0A0A",		-- 10, 10, 10, 10
        6674 => x"09090909",		-- 9, 9, 9, 9
        6675 => x"00000000",		-- 8, 8, 8, 8
        6676 => x"000B0A0B",		-- 8, 11, 10, 11
        6677 => x"0B0B0909",		-- 11, 11, 9, 9
        6678 => x"09090909",		-- 9, 9, 9, 9
        6679 => x"090B0000",		-- 9, 11, 8, 8
        6680 => x"000B0A0B",		-- 8, 11, 10, 11
        6681 => x"0B090909",		-- 11, 9, 9, 9
        6682 => x"0A0A0A09",		-- 10, 10, 10, 9
        6683 => x"0B0B0B00",		-- 11, 11, 11, 8
        6684 => x"000B000B",		-- 8, 11, 8, 11
        6685 => x"0B090909",		-- 11, 9, 9, 9
        6686 => x"0A0A0A0B",		-- 10, 10, 10, 11
        6687 => x"0B0B0B00",		-- 11, 11, 11, 8
        6688 => x"000B0000",		-- 8, 11, 8, 8
        6689 => x"000B0909",		-- 8, 11, 9, 9
        6690 => x"090A0A0B",		-- 9, 10, 10, 11
        6691 => x"0B0B0B00",		-- 11, 11, 11, 8
        6692 => x"000B0000",		-- 8, 11, 8, 8
        6693 => x"000B0B0B",		-- 8, 11, 11, 11
        6694 => x"0B09090B",		-- 11, 9, 9, 11
        6695 => x"0B090000",		-- 11, 9, 8, 8
        6696 => x"00000000",		-- 8, 8, 8, 8
        6697 => x"00090909",		-- 8, 9, 9, 9
        6698 => x"09090909",		-- 9, 9, 9, 9
        6699 => x"09090900",		-- 9, 9, 9, 8
        6700 => x"00000000",		-- 8, 8, 8, 8
        6701 => x"00000000",		-- 8, 8, 8, 8
        6702 => x"0B0B0B0B",		-- 11, 11, 11, 11
        6703 => x"00000000",		-- 8, 8, 8, 8
        6704 => x"00000000",		-- 8, 8, 8, 8
        6705 => x"0000000B",		-- 8, 8, 8, 11
        6706 => x"0B0B0B0B",		-- 11, 11, 11, 11
        6707 => x"00000000",		-- 8, 8, 8, 8

                --  sprite 24
        6708 => x"00000000",		-- 8, 8, 8, 8
        6709 => x"00000000",		-- 8, 8, 8, 8
        6710 => x"00000000",		-- 8, 8, 8, 8
        6711 => x"00000000",		-- 8, 8, 8, 8
        6712 => x"00000000",		-- 8, 8, 8, 8
        6713 => x"00000009",		-- 8, 8, 8, 9
        6714 => x"09090900",		-- 9, 9, 9, 8
        6715 => x"00000000",		-- 8, 8, 8, 8
        6716 => x"00000000",		-- 8, 8, 8, 8
        6717 => x"0B0B0B0B",		-- 11, 11, 11, 11
        6718 => x"09090909",		-- 9, 9, 9, 9
        6719 => x"09000000",		-- 9, 8, 8, 8
        6720 => x"0000000B",		-- 8, 8, 8, 11
        6721 => x"0B0B0B0B",		-- 11, 11, 11, 11
        6722 => x"0B09090A",		-- 11, 9, 9, 10
        6723 => x"09090900",		-- 9, 9, 9, 8
        6724 => x"000B0B00",		-- 8, 11, 11, 8
        6725 => x"0B0B0B0B",		-- 11, 11, 11, 11
        6726 => x"0B0B0A0A",		-- 11, 11, 10, 10
        6727 => x"09090909",		-- 9, 9, 9, 9
        6728 => x"000B0B00",		-- 8, 11, 11, 8
        6729 => x"0A090A0A",		-- 10, 9, 10, 10
        6730 => x"0B0A0A0A",		-- 11, 10, 10, 10
        6731 => x"09090009",		-- 9, 9, 8, 9
        6732 => x"000A0B0A",		-- 8, 10, 11, 10
        6733 => x"0A0B0A0A",		-- 10, 11, 10, 10
        6734 => x"0B0A0A0B",		-- 11, 10, 10, 11
        6735 => x"0B090000",		-- 11, 9, 8, 8
        6736 => x"000A0B00",		-- 8, 10, 11, 8
        6737 => x"0A0A0A0A",		-- 10, 10, 10, 10
        6738 => x"0A0A0B0B",		-- 10, 10, 11, 11
        6739 => x"0B000000",		-- 11, 8, 8, 8
        6740 => x"000A0B00",		-- 8, 10, 11, 8
        6741 => x"0A0A0A0A",		-- 10, 10, 10, 10
        6742 => x"09090909",		-- 9, 9, 9, 9
        6743 => x"00000000",		-- 8, 8, 8, 8
        6744 => x"000A0B0A",		-- 8, 10, 11, 10
        6745 => x"0B0B0A0A",		-- 11, 11, 10, 10
        6746 => x"0A09090B",		-- 10, 9, 9, 11
        6747 => x"0B090000",		-- 11, 9, 8, 8
        6748 => x"000A0B0A",		-- 8, 10, 11, 10
        6749 => x"0B090A0A",		-- 11, 9, 10, 10
        6750 => x"0A0B0B0B",		-- 10, 11, 11, 11
        6751 => x"0B0B0000",		-- 11, 11, 8, 8
        6752 => x"000A0B00",		-- 8, 10, 11, 8
        6753 => x"0B09090A",		-- 11, 9, 9, 10
        6754 => x"0A0B0B0B",		-- 10, 11, 11, 11
        6755 => x"0B0B0900",		-- 11, 11, 9, 8
        6756 => x"000A0B00",		-- 8, 10, 11, 8
        6757 => x"000B0909",		-- 8, 11, 9, 9
        6758 => x"090B0B0B",		-- 9, 11, 11, 11
        6759 => x"0B090900",		-- 11, 9, 9, 8
        6760 => x"000A0B00",		-- 8, 10, 11, 8
        6761 => x"090B0B0B",		-- 9, 11, 11, 11
        6762 => x"0B090909",		-- 11, 9, 9, 9
        6763 => x"09090B0B",		-- 9, 9, 11, 11
        6764 => x"000B0B0B",		-- 8, 11, 11, 11
        6765 => x"0B090909",		-- 11, 9, 9, 9
        6766 => x"09090909",		-- 9, 9, 9, 9
        6767 => x"090B0B0B",		-- 9, 11, 11, 11
        6768 => x"000B0B00",		-- 8, 11, 11, 8
        6769 => x"0B0B0B00",		-- 11, 11, 11, 8
        6770 => x"00000000",		-- 8, 8, 8, 8
        6771 => x"0B0B0B00",		-- 11, 11, 11, 8

                --  sprite 25
        6772 => x"00000000",		-- 8, 8, 8, 8
        6773 => x"00000009",		-- 8, 8, 8, 9
        6774 => x"09090900",		-- 9, 9, 9, 8
        6775 => x"00000000",		-- 8, 8, 8, 8
        6776 => x"00000000",		-- 8, 8, 8, 8
        6777 => x"0B0B0B0B",		-- 11, 11, 11, 11
        6778 => x"09090909",		-- 9, 9, 9, 9
        6779 => x"09000000",		-- 9, 8, 8, 8
        6780 => x"0000000B",		-- 8, 8, 8, 11
        6781 => x"0B0B0B0B",		-- 11, 11, 11, 11
        6782 => x"0B09090A",		-- 11, 9, 9, 10
        6783 => x"09090900",		-- 9, 9, 9, 8
        6784 => x"0B0B0000",		-- 11, 11, 8, 8
        6785 => x"0B0B0B0B",		-- 11, 11, 11, 11
        6786 => x"0B0B0A0A",		-- 11, 11, 10, 10
        6787 => x"09090909",		-- 9, 9, 9, 9
        6788 => x"0B0B0000",		-- 11, 11, 8, 8
        6789 => x"0A090A0A",		-- 10, 9, 10, 10
        6790 => x"0B0A0A0A",		-- 11, 10, 10, 10
        6791 => x"09090009",		-- 9, 9, 8, 9
        6792 => x"0A0B0A0A",		-- 10, 11, 10, 10
        6793 => x"0A0B0A0A",		-- 10, 11, 10, 10
        6794 => x"0B0A0A0B",		-- 11, 10, 10, 11
        6795 => x"0B090000",		-- 11, 9, 8, 8
        6796 => x"0A0B0000",		-- 10, 11, 8, 8
        6797 => x"0A0A0A0A",		-- 10, 10, 10, 10
        6798 => x"0A0A0B0B",		-- 10, 10, 11, 11
        6799 => x"0B000000",		-- 11, 8, 8, 8
        6800 => x"0A0B0000",		-- 10, 11, 8, 8
        6801 => x"0A0A0A0A",		-- 10, 10, 10, 10
        6802 => x"09090909",		-- 9, 9, 9, 9
        6803 => x"00000000",		-- 8, 8, 8, 8
        6804 => x"0A0B0A0B",		-- 10, 11, 10, 11
        6805 => x"0B0B0909",		-- 11, 11, 9, 9
        6806 => x"09090909",		-- 9, 9, 9, 9
        6807 => x"090B0000",		-- 9, 11, 8, 8
        6808 => x"0A0B0A0B",		-- 10, 11, 10, 11
        6809 => x"0B090909",		-- 11, 9, 9, 9
        6810 => x"0A0A0A09",		-- 10, 10, 10, 9
        6811 => x"0B0B0B00",		-- 11, 11, 11, 8
        6812 => x"0A0B000B",		-- 10, 11, 8, 11
        6813 => x"0B090909",		-- 11, 9, 9, 9
        6814 => x"0A0A0A0B",		-- 10, 10, 10, 11
        6815 => x"0B0B0B00",		-- 11, 11, 11, 8
        6816 => x"0A0B0000",		-- 10, 11, 8, 8
        6817 => x"000B0909",		-- 8, 11, 9, 9
        6818 => x"090A0A0B",		-- 9, 10, 10, 11
        6819 => x"0B0B0B00",		-- 11, 11, 11, 8
        6820 => x"0A0B0000",		-- 10, 11, 8, 8
        6821 => x"000B0B0B",		-- 8, 11, 11, 11
        6822 => x"0B09090B",		-- 11, 9, 9, 11
        6823 => x"0B090000",		-- 11, 9, 8, 8
        6824 => x"0B0B0000",		-- 11, 11, 8, 8
        6825 => x"00090909",		-- 8, 9, 9, 9
        6826 => x"09090909",		-- 9, 9, 9, 9
        6827 => x"09090900",		-- 9, 9, 9, 8
        6828 => x"0B0B0000",		-- 11, 11, 8, 8
        6829 => x"00000000",		-- 8, 8, 8, 8
        6830 => x"0B0B0B0B",		-- 11, 11, 11, 11
        6831 => x"00000000",		-- 8, 8, 8, 8
        6832 => x"00000000",		-- 8, 8, 8, 8
        6833 => x"0000000B",		-- 8, 8, 8, 11
        6834 => x"0B0B0B0B",		-- 11, 11, 11, 11
        6835 => x"00000000",		-- 8, 8, 8, 8

                --  sprite 26
        6836 => x"00000000",		-- 8, 8, 8, 8
        6837 => x"00000000",		-- 8, 8, 8, 8
        6838 => x"00000000",		-- 8, 8, 8, 8
        6839 => x"00000000",		-- 8, 8, 8, 8
        6840 => x"00000000",		-- 8, 8, 8, 8
        6841 => x"00000909",		-- 8, 8, 9, 9
        6842 => x"09090000",		-- 9, 9, 8, 8
        6843 => x"00000000",		-- 8, 8, 8, 8
        6844 => x"0000000B",		-- 8, 8, 8, 11
        6845 => x"0B0B0B09",		-- 11, 11, 11, 9
        6846 => x"09090909",		-- 9, 9, 9, 9
        6847 => x"00000000",		-- 8, 8, 8, 8
        6848 => x"00000B0B",		-- 8, 8, 11, 11
        6849 => x"0B0B0B0B",		-- 11, 11, 11, 11
        6850 => x"09090A09",		-- 9, 9, 10, 9
        6851 => x"09000000",		-- 9, 8, 8, 8
        6852 => x"0000000B",		-- 8, 8, 8, 11
        6853 => x"0B0B0B0B",		-- 11, 11, 11, 11
        6854 => x"0B0A0A09",		-- 11, 10, 10, 9
        6855 => x"09000000",		-- 9, 8, 8, 8
        6856 => x"0000000A",		-- 8, 8, 8, 10
        6857 => x"090A0A0B",		-- 9, 10, 10, 11
        6858 => x"0A0A0A09",		-- 10, 10, 10, 9
        6859 => x"09090000",		-- 9, 9, 8, 8
        6860 => x"000A0A0A",		-- 8, 10, 10, 10
        6861 => x"0B0A0A0B",		-- 11, 10, 10, 11
        6862 => x"0A0A0B0B",		-- 10, 10, 11, 11
        6863 => x"09090900",		-- 9, 9, 9, 8
        6864 => x"0000000A",		-- 8, 8, 8, 10
        6865 => x"0A0A0A0A",		-- 10, 10, 10, 10
        6866 => x"0A0B0B0B",		-- 10, 11, 11, 11
        6867 => x"00000900",		-- 8, 8, 9, 8
        6868 => x"00000A0A",		-- 8, 8, 10, 10
        6869 => x"0A0A0A09",		-- 10, 10, 10, 9
        6870 => x"09090909",		-- 9, 9, 9, 9
        6871 => x"00000000",		-- 8, 8, 8, 8
        6872 => x"00000A0A",		-- 8, 8, 10, 10
        6873 => x"0A0B0B0B",		-- 10, 11, 11, 11
        6874 => x"0B0B0B09",		-- 11, 11, 11, 9
        6875 => x"09000000",		-- 9, 8, 8, 8
        6876 => x"0000000A",		-- 8, 8, 8, 10
        6877 => x"0A0B0B0B",		-- 10, 11, 11, 11
        6878 => x"0B0B0B0B",		-- 11, 11, 11, 11
        6879 => x"09000000",		-- 9, 8, 8, 8
        6880 => x"00000000",		-- 8, 8, 8, 8
        6881 => x"090B0B0B",		-- 9, 11, 11, 11
        6882 => x"0B0B0B0B",		-- 11, 11, 11, 11
        6883 => x"09090000",		-- 9, 9, 8, 8
        6884 => x"0000000B",		-- 8, 8, 8, 11
        6885 => x"0B090909",		-- 11, 9, 9, 9
        6886 => x"0B0B0B09",		-- 11, 11, 11, 9
        6887 => x"09090900",		-- 9, 9, 9, 8
        6888 => x"0000000B",		-- 8, 8, 8, 11
        6889 => x"0B0B0B0B",		-- 11, 11, 11, 11
        6890 => x"09090909",		-- 9, 9, 9, 9
        6891 => x"09090B0B",		-- 9, 9, 11, 11
        6892 => x"00000B0B",		-- 8, 8, 11, 11
        6893 => x"09090909",		-- 9, 9, 9, 9
        6894 => x"09090909",		-- 9, 9, 9, 9
        6895 => x"090B0B0B",		-- 9, 11, 11, 11
        6896 => x"000B0B0B",		-- 8, 11, 11, 11
        6897 => x"0B000000",		-- 11, 8, 8, 8
        6898 => x"00000000",		-- 8, 8, 8, 8
        6899 => x"0B0B0B00",		-- 11, 11, 11, 8

--		****  MAP  ****
        6900 => x"00000016", -- pedding 
        6901 => x"00000016", -- pedding 
        6902 => x"00000016", -- pedding 
        6903 => x"00000016", -- pedding 
        6904 => x"00000016", -- pedding 
        6905 => x"00000016", -- pedding 
        6906 => x"00000016", -- pedding 
        6907 => x"00000016", -- pedding 
        6908 => x"00000016", -- pedding 
        6909 => x"00000016", -- pedding 
        6910 => x"00000016", -- pedding 
        6911 => x"00000016", -- pedding 
        6912 => x"00000016", -- pedding 
        6913 => x"00000016", -- pedding 
        6914 => x"00000016", -- pedding 
        6915 => x"00000016", -- pedding 
        6916 => x"00000016", -- pedding 
        6917 => x"00000016", -- pedding 
        6918 => x"00000016", -- pedding 
        6919 => x"00000016", -- pedding 
        6920 => x"00000016", -- pedding 
        6921 => x"00000016", -- pedding 
        6922 => x"00000016", -- pedding 
        6923 => x"00000016", -- pedding 
        6924 => x"00000016", -- pedding 
        6925 => x"00000016", -- pedding 
        6926 => x"00000016", -- pedding 
        6927 => x"00000016", -- pedding 
        6928 => x"00000016", -- pedding 
        6929 => x"00000016", -- pedding 
        6930 => x"00000016", -- pedding 
        6931 => x"00000016", -- pedding 
        6932 => x"00000016", -- pedding 
        6933 => x"00000016", -- pedding 
        6934 => x"00000016", -- pedding 
        6935 => x"00000016", -- pedding 
        6936 => x"00000016", -- pedding 
        6937 => x"00000016", -- pedding 
        6938 => x"00000016", -- pedding 
        6939 => x"00000016", -- pedding 
        6940 => x"00000016", -- pedding 
        6941 => x"00000016", -- pedding 
        6942 => x"00000016", -- pedding 
        6943 => x"00000016", -- pedding 
        6944 => x"00000016", -- pedding 
        6945 => x"00000016", -- pedding 
        6946 => x"00000016", -- pedding 
        6947 => x"00000016", -- pedding 
        6948 => x"00000016", -- pedding 
        6949 => x"00000016", -- pedding 
        6950 => x"00000016", -- pedding 
        6951 => x"00000016", -- pedding 
        6952 => x"00000016", -- pedding 
        6953 => x"00000016", -- pedding 
        6954 => x"00000016", -- pedding 
        6955 => x"00000016", -- pedding 
        6956 => x"00000016", -- pedding 
        6957 => x"00000016", -- pedding 
        6958 => x"00000016", -- pedding 
        6959 => x"00000016", -- pedding 
        6960 => x"00000016", -- pedding 
        6961 => x"00000016", -- pedding 
        6962 => x"00000016", -- pedding 
        6963 => x"00000016", -- pedding 
        6964 => x"00000016", -- pedding 
        6965 => x"00000016", -- pedding 
        6966 => x"00000016", -- pedding 
        6967 => x"00000016", -- pedding 
        6968 => x"00000016", -- pedding 
        6969 => x"00000016", -- pedding 
        6970 => x"00000016", -- pedding 
        6971 => x"00000016", -- pedding 
        6972 => x"00000016", -- pedding 
        6973 => x"00000016", -- pedding 
        6974 => x"00000016", -- pedding 
        6975 => x"00000016", -- pedding 
        6976 => x"00000016", -- pedding 
        6977 => x"00000016", -- pedding 
        6978 => x"00000016", -- pedding 
        6979 => x"00000016", -- pedding 
        6980 => x"00000016", -- pedding 
        6981 => x"00000016", -- pedding 
        6982 => x"00000016", -- pedding 
        6983 => x"00000016", -- pedding 
        6984 => x"00000016", -- pedding 
        6985 => x"00000016", -- pedding 
        6986 => x"00000016", -- pedding 
        6987 => x"00000016", -- pedding 
        6988 => x"00000016", -- pedding 
        6989 => x"00000016", -- pedding 
        6990 => x"00000016", -- pedding 
        6991 => x"00000016", -- pedding 
        6992 => x"00000016", -- pedding 
        6993 => x"00000016", -- pedding 
        6994 => x"00000016", -- pedding 
        6995 => x"00000016", -- pedding 
        6996 => x"00000016", -- pedding 
        6997 => x"00000016", -- pedding 
        6998 => x"00000016", -- pedding 
        6999 => x"00000016", -- pedding 
        7000 => x"00000016", -- pedding 
        7001 => x"00000016", -- pedding 
        7002 => x"00000016", -- pedding 
        7003 => x"00000016", -- pedding 
        7004 => x"00000016", -- pedding 
        7005 => x"00000016", -- pedding 
        7006 => x"00000016", -- pedding 
        7007 => x"00000016", -- pedding 
        7008 => x"00000016", -- pedding 
        7009 => x"00000016", -- pedding 
        7010 => x"00000016", -- pedding 
        7011 => x"00000016", -- pedding 
        7012 => x"00000016", -- pedding 
        7013 => x"00000016", -- pedding 
        7014 => x"00000016", -- pedding 
        7015 => x"00000016", -- pedding 
        7016 => x"00000016", -- pedding 
        7017 => x"00000016", -- pedding 
        7018 => x"00000016", -- pedding 
        7019 => x"00000016", -- pedding 
        7020 => x"00000016", -- pedding 
        7021 => x"00000016", -- pedding 
        7022 => x"00000016", -- pedding 
        7023 => x"00000016", -- pedding 
        7024 => x"00000016", -- pedding 
        7025 => x"00000016", -- pedding 
        7026 => x"00000016", -- pedding 
        7027 => x"00000016", -- pedding 
        7028 => x"00000016", -- pedding 
        7029 => x"00000016", -- pedding 
        7030 => x"00000016", -- pedding 
        7031 => x"00000016", -- pedding 
        7032 => x"00000016", -- header 
        7033 => x"00000016", -- header 
        7034 => x"00000016", -- header 
        7035 => x"00000016", -- header 
        7036 => x"00000016", -- header 
        7037 => x"00000016", -- header 
        7038 => x"00000016", -- header 
        7039 => x"00000016", -- header 
        7040 => x"00000016", -- header 
        7041 => x"00000016", -- header 
        7042 => x"00000016", -- header 
        7043 => x"00000016", -- header 
        7044 => x"00000016", -- header 
        7045 => x"00000016", -- header 
        7046 => x"00000016", -- header 
        7047 => x"00000016", -- header 
        7048 => x"00000016", -- pedding 
        7049 => x"00000016", -- pedding 
        7050 => x"00000016", -- pedding 
        7051 => x"00000016", -- pedding 
        7052 => x"00000016", -- pedding 
        7053 => x"00000016", -- pedding 
        7054 => x"00000016", -- pedding 
        7055 => x"00000016", -- pedding 
        7056 => x"00000016", -- pedding 
        7057 => x"00000016", -- pedding 
        7058 => x"00000016", -- pedding 
        7059 => x"00000016", -- pedding 
        7060 => x"00000016", -- pedding 
        7061 => x"00000016", -- pedding 
        7062 => x"00000016", -- pedding 
        7063 => x"00000016", -- pedding 
        7064 => x"00000016", -- pedding 
        7065 => x"00000016", -- pedding 
        7066 => x"00000016", -- pedding 
        7067 => x"00000016", -- pedding 
        7068 => x"00000016", -- pedding 
        7069 => x"00000016", -- pedding 
        7070 => x"00000016", -- pedding 
        7071 => x"00000016", -- pedding 
        7072 => x"00000016", -- header 
        7073 => x"00000016", -- header 
        7074 => x"00000016", -- header 
        7075 => x"00000016", -- header 
        7076 => x"00000016", -- header 
        7077 => x"00000016", -- header 
        7078 => x"00000016", -- header 
        7079 => x"00000016", -- header 
        7080 => x"00000016", -- header 
        7081 => x"00000016", -- header 
        7082 => x"00000016", -- header 
        7083 => x"00000016", -- header 
        7084 => x"00000016", -- header 
        7085 => x"00000016", -- header 
        7086 => x"00000016", -- header 
        7087 => x"00000016", -- header 
        7088 => x"00000016", -- pedding 
        7089 => x"00000016", -- pedding 
        7090 => x"00000016", -- pedding 
        7091 => x"00000016", -- pedding 
        7092 => x"00000016", -- pedding 
        7093 => x"00000016", -- pedding 
        7094 => x"00000016", -- pedding 
        7095 => x"00000016", -- pedding 
        7096 => x"00000016", -- pedding 
        7097 => x"00000016", -- pedding 
        7098 => x"00000016", -- pedding 
        7099 => x"00000016", -- pedding 
        7100 => x"00000016", -- pedding 
        7101 => x"00000016", -- pedding 
        7102 => x"00000016", -- pedding 
        7103 => x"00000016", -- pedding 
        7104 => x"00000016", -- pedding 
        7105 => x"00000016", -- pedding 
        7106 => x"00000016", -- pedding 
        7107 => x"00000016", -- pedding 
        7108 => x"00000016", -- pedding 
        7109 => x"00000016", -- pedding 
        7110 => x"00000016", -- pedding 
        7111 => x"00000016", -- pedding 
        7112 => x"00000016", -- header 
        7113 => x"00000016", -- header 
        7114 => x"00000016", -- header 
        7115 => x"00000016", -- header 
        7116 => x"00000016", -- header 
        7117 => x"00000016", -- header 
        7118 => x"00000016", -- header 
        7119 => x"00000016", -- header 
        7120 => x"00000016", -- header 
        7121 => x"00000016", -- header 
        7122 => x"00000016", -- header 
        7123 => x"00000016", -- header 
        7124 => x"00000016", -- header 
        7125 => x"00000016", -- header 
        7126 => x"00000016", -- header 
        7127 => x"00000016", -- header 
        7128 => x"00000016", -- pedding 
        7129 => x"00000016", -- pedding 
        7130 => x"00000016", -- pedding 
        7131 => x"00000016", -- pedding 
        7132 => x"00000016", -- pedding 
        7133 => x"00000016", -- pedding 
        7134 => x"00000016", -- pedding 
        7135 => x"00000016", -- pedding 
        7136 => x"00000016", -- pedding 
        7137 => x"00000016", -- pedding 
        7138 => x"00000016", -- pedding 
        7139 => x"00000016", -- pedding 
        7140 => x"00000016", -- pedding 
        7141 => x"00000016", -- pedding 
        7142 => x"00000016", -- pedding 
        7143 => x"00000016", -- pedding 
        7144 => x"00000016", -- pedding 
        7145 => x"00000016", -- pedding 
        7146 => x"00000016", -- pedding 
        7147 => x"00000016", -- pedding 
        7148 => x"00000016", -- pedding 
        7149 => x"00000016", -- pedding 
        7150 => x"00000016", -- pedding 
        7151 => x"00000016", -- pedding 
        7152 => x"00000016", -- header 
        7153 => x"00000016", -- header 
        7154 => x"00000016", -- header 
        7155 => x"00000016", -- header 
        7156 => x"00000016", -- header 
        7157 => x"00000016", -- header 
        7158 => x"00000016", -- header 
        7159 => x"00000016", -- header 
        7160 => x"00000016", -- header 
        7161 => x"00000016", -- header 
        7162 => x"00000016", -- header 
        7163 => x"00000016", -- header 
        7164 => x"00000016", -- header 
        7165 => x"00000016", -- header 
        7166 => x"00000016", -- header 
        7167 => x"00000016", -- header 
        7168 => x"00000016", -- pedding 
        7169 => x"00000016", -- pedding 
        7170 => x"00000016", -- pedding 
        7171 => x"00000016", -- pedding 
        7172 => x"00000016", -- pedding 
        7173 => x"00000016", -- pedding 
        7174 => x"00000016", -- pedding 
        7175 => x"00000016", -- pedding 
        7176 => x"00000016", -- pedding 
        7177 => x"00000016", -- pedding 
        7178 => x"00000016", -- pedding 
        7179 => x"00000016", -- pedding 
        7180 => x"00000016", -- pedding 
        7181 => x"00000016", -- pedding 
        7182 => x"00000016", -- pedding 
        7183 => x"00000016", -- pedding 
        7184 => x"00000016", -- pedding 
        7185 => x"00000016", -- pedding 
        7186 => x"00000016", -- pedding 
        7187 => x"00000016", -- pedding 
        7188 => x"00000016", -- pedding 
        7189 => x"00000016", -- pedding 
        7190 => x"00000016", -- pedding 
        7191 => x"00000016", -- pedding 
        7192 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7193 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7194 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7195 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7196 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7197 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7198 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7199 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7200 => x"00000001", -- z: 0 rot: 0 ptr: 319
        7201 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7202 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7203 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7204 => x"00000001", -- z: 0 rot: 0 ptr: 319
        7205 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7206 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7207 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7208 => x"00000016", -- pedding 
        7209 => x"00000016", -- pedding 
        7210 => x"00000016", -- pedding 
        7211 => x"00000016", -- pedding 
        7212 => x"00000016", -- pedding 
        7213 => x"00000016", -- pedding 
        7214 => x"00000016", -- pedding 
        7215 => x"00000016", -- pedding 
        7216 => x"00000016", -- pedding 
        7217 => x"00000016", -- pedding 
        7218 => x"00000016", -- pedding 
        7219 => x"00000016", -- pedding 
        7220 => x"00000016", -- pedding 
        7221 => x"00000016", -- pedding 
        7222 => x"00000016", -- pedding 
        7223 => x"00000016", -- pedding 
        7224 => x"00000016", -- pedding 
        7225 => x"00000016", -- pedding 
        7226 => x"00000016", -- pedding 
        7227 => x"00000016", -- pedding 
        7228 => x"00000016", -- pedding 
        7229 => x"00000016", -- pedding 
        7230 => x"00000016", -- pedding 
        7231 => x"00000016", -- pedding 
        7232 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7233 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7234 => x"00000003", -- z: 0 rot: 0 ptr: 447
        7235 => x"00000005", -- z: 0 rot: 0 ptr: 575
        7236 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7237 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7238 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7239 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7240 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7241 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7242 => x"00000001", -- z: 0 rot: 0 ptr: 319
        7243 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7244 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7245 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7246 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7247 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7248 => x"00000016", -- pedding 
        7249 => x"00000016", -- pedding 
        7250 => x"00000016", -- pedding 
        7251 => x"00000016", -- pedding 
        7252 => x"00000016", -- pedding 
        7253 => x"00000016", -- pedding 
        7254 => x"00000016", -- pedding 
        7255 => x"00000016", -- pedding 
        7256 => x"00000016", -- pedding 
        7257 => x"00000016", -- pedding 
        7258 => x"00000016", -- pedding 
        7259 => x"00000016", -- pedding 
        7260 => x"00000016", -- pedding 
        7261 => x"00000016", -- pedding 
        7262 => x"00000016", -- pedding 
        7263 => x"00000016", -- pedding 
        7264 => x"00000016", -- pedding 
        7265 => x"00000016", -- pedding 
        7266 => x"00000016", -- pedding 
        7267 => x"00000016", -- pedding 
        7268 => x"00000016", -- pedding 
        7269 => x"00000016", -- pedding 
        7270 => x"00000016", -- pedding 
        7271 => x"00000016", -- pedding 
        7272 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7273 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7274 => x"00000015", -- z: 0 rot: 0 ptr: 831
        7275 => x"00000017", -- z: 0 rot: 0 ptr: 959
        7276 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7277 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7278 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7279 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7280 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7281 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7282 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7283 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7284 => x"00000001", -- z: 0 rot: 0 ptr: 319
        7285 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7286 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7287 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7288 => x"00000016", -- pedding 
        7289 => x"00000016", -- pedding 
        7290 => x"00000016", -- pedding 
        7291 => x"00000016", -- pedding 
        7292 => x"00000016", -- pedding 
        7293 => x"00000016", -- pedding 
        7294 => x"00000016", -- pedding 
        7295 => x"00000016", -- pedding 
        7296 => x"00000016", -- pedding 
        7297 => x"00000016", -- pedding 
        7298 => x"00000016", -- pedding 
        7299 => x"00000016", -- pedding 
        7300 => x"00000016", -- pedding 
        7301 => x"00000016", -- pedding 
        7302 => x"00000016", -- pedding 
        7303 => x"00000016", -- pedding 
        7304 => x"00000016", -- pedding 
        7305 => x"00000016", -- pedding 
        7306 => x"00000016", -- pedding 
        7307 => x"00000016", -- pedding 
        7308 => x"00000016", -- pedding 
        7309 => x"00000016", -- pedding 
        7310 => x"00000016", -- pedding 
        7311 => x"00000016", -- pedding 
        7312 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7313 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7314 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7315 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7316 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7317 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7318 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7319 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7320 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7321 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7322 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7323 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7324 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7325 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7326 => x"00000024", -- z: 0 rot: 0 ptr: 1023
        7327 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7328 => x"00000016", -- pedding 
        7329 => x"00000016", -- pedding 
        7330 => x"00000016", -- pedding 
        7331 => x"00000016", -- pedding 
        7332 => x"00000016", -- pedding 
        7333 => x"00000016", -- pedding 
        7334 => x"00000016", -- pedding 
        7335 => x"00000016", -- pedding 
        7336 => x"00000016", -- pedding 
        7337 => x"00000016", -- pedding 
        7338 => x"00000016", -- pedding 
        7339 => x"00000016", -- pedding 
        7340 => x"00000016", -- pedding 
        7341 => x"00000016", -- pedding 
        7342 => x"00000016", -- pedding 
        7343 => x"00000016", -- pedding 
        7344 => x"00000016", -- pedding 
        7345 => x"00000016", -- pedding 
        7346 => x"00000016", -- pedding 
        7347 => x"00000016", -- pedding 
        7348 => x"00000016", -- pedding 
        7349 => x"00000016", -- pedding 
        7350 => x"00000016", -- pedding 
        7351 => x"00000016", -- pedding 
        7352 => x"00000025", -- z: 0 rot: 0 ptr: 1087
        7353 => x"00000025", -- z: 0 rot: 0 ptr: 1087
        7354 => x"00000025", -- z: 0 rot: 0 ptr: 1087
        7355 => x"00000025", -- z: 0 rot: 0 ptr: 1087
        7356 => x"00000025", -- z: 0 rot: 0 ptr: 1087
        7357 => x"00000025", -- z: 0 rot: 0 ptr: 1087
        7358 => x"00000025", -- z: 0 rot: 0 ptr: 1087
        7359 => x"00000025", -- z: 0 rot: 0 ptr: 1087
        7360 => x"00000025", -- z: 0 rot: 0 ptr: 1087
        7361 => x"00000025", -- z: 0 rot: 0 ptr: 1087
        7362 => x"00000025", -- z: 0 rot: 0 ptr: 1087
        7363 => x"00000025", -- z: 0 rot: 0 ptr: 1087
        7364 => x"00000025", -- z: 0 rot: 0 ptr: 1087
        7365 => x"00000025", -- z: 0 rot: 0 ptr: 1087
        7366 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7367 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7368 => x"00000016", -- pedding 
        7369 => x"00000016", -- pedding 
        7370 => x"00000016", -- pedding 
        7371 => x"00000016", -- pedding 
        7372 => x"00000016", -- pedding 
        7373 => x"00000016", -- pedding 
        7374 => x"00000016", -- pedding 
        7375 => x"00000016", -- pedding 
        7376 => x"00000016", -- pedding 
        7377 => x"00000016", -- pedding 
        7378 => x"00000016", -- pedding 
        7379 => x"00000016", -- pedding 
        7380 => x"00000016", -- pedding 
        7381 => x"00000016", -- pedding 
        7382 => x"00000016", -- pedding 
        7383 => x"00000016", -- pedding 
        7384 => x"00000016", -- pedding 
        7385 => x"00000016", -- pedding 
        7386 => x"00000016", -- pedding 
        7387 => x"00000016", -- pedding 
        7388 => x"00000016", -- pedding 
        7389 => x"00000016", -- pedding 
        7390 => x"00000016", -- pedding 
        7391 => x"00000016", -- pedding 
        7392 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7393 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7394 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7395 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7396 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7397 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7398 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7399 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7400 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7401 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7402 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7403 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7404 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7405 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7406 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7407 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7408 => x"00000016", -- pedding 
        7409 => x"00000016", -- pedding 
        7410 => x"00000016", -- pedding 
        7411 => x"00000016", -- pedding 
        7412 => x"00000016", -- pedding 
        7413 => x"00000016", -- pedding 
        7414 => x"00000016", -- pedding 
        7415 => x"00000016", -- pedding 
        7416 => x"00000016", -- pedding 
        7417 => x"00000016", -- pedding 
        7418 => x"00000016", -- pedding 
        7419 => x"00000016", -- pedding 
        7420 => x"00000016", -- pedding 
        7421 => x"00000016", -- pedding 
        7422 => x"00000016", -- pedding 
        7423 => x"00000016", -- pedding 
        7424 => x"00000016", -- pedding 
        7425 => x"00000016", -- pedding 
        7426 => x"00000016", -- pedding 
        7427 => x"00000016", -- pedding 
        7428 => x"00000016", -- pedding 
        7429 => x"00000016", -- pedding 
        7430 => x"00000016", -- pedding 
        7431 => x"00000016", -- pedding 
        7432 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7433 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7434 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7435 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7436 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7437 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7438 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7439 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7440 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7441 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7442 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7443 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7444 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7445 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7446 => x"00000013", -- z: 0 rot: 0 ptr: 703
        7447 => x"00000013", -- z: 0 rot: 0 ptr: 703
        7448 => x"00000016", -- pedding 
        7449 => x"00000016", -- pedding 
        7450 => x"00000016", -- pedding 
        7451 => x"00000016", -- pedding 
        7452 => x"00000016", -- pedding 
        7453 => x"00000016", -- pedding 
        7454 => x"00000016", -- pedding 
        7455 => x"00000016", -- pedding 
        7456 => x"00000016", -- pedding 
        7457 => x"00000016", -- pedding 
        7458 => x"00000016", -- pedding 
        7459 => x"00000016", -- pedding 
        7460 => x"00000016", -- pedding 
        7461 => x"00000016", -- pedding 
        7462 => x"00000016", -- pedding 
        7463 => x"00000016", -- pedding 
        7464 => x"00000016", -- pedding 
        7465 => x"00000016", -- pedding 
        7466 => x"00000016", -- pedding 
        7467 => x"00000016", -- pedding 
        7468 => x"00000016", -- pedding 
        7469 => x"00000016", -- pedding 
        7470 => x"00000016", -- pedding 
        7471 => x"00000016", -- pedding 
        7472 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7473 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7474 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7475 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7476 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7477 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7478 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7479 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7480 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7481 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7482 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7483 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7484 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7485 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7486 => x"00000013", -- z: 0 rot: 0 ptr: 703
        7487 => x"00000013", -- z: 0 rot: 0 ptr: 703
        7488 => x"00000016", -- pedding 
        7489 => x"00000016", -- pedding 
        7490 => x"00000016", -- pedding 
        7491 => x"00000016", -- pedding 
        7492 => x"00000016", -- pedding 
        7493 => x"00000016", -- pedding 
        7494 => x"00000016", -- pedding 
        7495 => x"00000016", -- pedding 
        7496 => x"00000016", -- pedding 
        7497 => x"00000016", -- pedding 
        7498 => x"00000016", -- pedding 
        7499 => x"00000016", -- pedding 
        7500 => x"00000016", -- pedding 
        7501 => x"00000016", -- pedding 
        7502 => x"00000016", -- pedding 
        7503 => x"00000016", -- pedding 
        7504 => x"00000016", -- pedding 
        7505 => x"00000016", -- pedding 
        7506 => x"00000016", -- pedding 
        7507 => x"00000016", -- pedding 
        7508 => x"00000016", -- pedding 
        7509 => x"00000016", -- pedding 
        7510 => x"00000016", -- pedding 
        7511 => x"00000016", -- pedding 
        7512 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7513 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7514 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7515 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7516 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7517 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7518 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7519 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7520 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7521 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7522 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7523 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7524 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7525 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7526 => x"00000013", -- z: 0 rot: 0 ptr: 703
        7527 => x"00000013", -- z: 0 rot: 0 ptr: 703
        7528 => x"00000016", -- pedding 
        7529 => x"00000016", -- pedding 
        7530 => x"00000016", -- pedding 
        7531 => x"00000016", -- pedding 
        7532 => x"00000016", -- pedding 
        7533 => x"00000016", -- pedding 
        7534 => x"00000016", -- pedding 
        7535 => x"00000016", -- pedding 
        7536 => x"00000016", -- pedding 
        7537 => x"00000016", -- pedding 
        7538 => x"00000016", -- pedding 
        7539 => x"00000016", -- pedding 
        7540 => x"00000016", -- pedding 
        7541 => x"00000016", -- pedding 
        7542 => x"00000016", -- pedding 
        7543 => x"00000016", -- pedding 
        7544 => x"00000016", -- pedding 
        7545 => x"00000016", -- pedding 
        7546 => x"00000016", -- pedding 
        7547 => x"00000016", -- pedding 
        7548 => x"00000016", -- pedding 
        7549 => x"00000016", -- pedding 
        7550 => x"00000016", -- pedding 
        7551 => x"00000016", -- pedding 
        7552 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7553 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7554 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7555 => x"00000092", -- z: 0 rot: 0 ptr: 3455
        7556 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7557 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7558 => x"00000092", -- z: 0 rot: 0 ptr: 3455
        7559 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7560 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7561 => x"00000092", -- z: 0 rot: 0 ptr: 3455
        7562 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7563 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7564 => x"00000092", -- z: 0 rot: 0 ptr: 3455
        7565 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7566 => x"00000013", -- z: 0 rot: 0 ptr: 703
        7567 => x"00000013", -- z: 0 rot: 0 ptr: 703
        7568 => x"00000016", -- pedding 
        7569 => x"00000016", -- pedding 
        7570 => x"00000016", -- pedding 
        7571 => x"00000016", -- pedding 
        7572 => x"00000016", -- pedding 
        7573 => x"00000016", -- pedding 
        7574 => x"00000016", -- pedding 
        7575 => x"00000016", -- pedding 
        7576 => x"00000016", -- pedding 
        7577 => x"00000016", -- pedding 
        7578 => x"00000016", -- pedding 
        7579 => x"00000016", -- pedding 
        7580 => x"00000016", -- pedding 
        7581 => x"00000016", -- pedding 
        7582 => x"00000016", -- pedding 
        7583 => x"00000016", -- pedding 
        7584 => x"00000016", -- pedding 
        7585 => x"00000016", -- pedding 
        7586 => x"00000016", -- pedding 
        7587 => x"00000016", -- pedding 
        7588 => x"00000016", -- pedding 
        7589 => x"00000016", -- pedding 
        7590 => x"00000016", -- pedding 
        7591 => x"00000016", -- pedding 
        7592 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7593 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7594 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7595 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7596 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7597 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7598 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7599 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7600 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7601 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7602 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7603 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7604 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7605 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7606 => x"00000013", -- z: 0 rot: 0 ptr: 703
        7607 => x"00000013", -- z: 0 rot: 0 ptr: 703
        7608 => x"00000016", -- pedding 
        7609 => x"00000016", -- pedding 
        7610 => x"00000016", -- pedding 
        7611 => x"00000016", -- pedding 
        7612 => x"00000016", -- pedding 
        7613 => x"00000016", -- pedding 
        7614 => x"00000016", -- pedding 
        7615 => x"00000016", -- pedding 
        7616 => x"00000016", -- pedding 
        7617 => x"00000016", -- pedding 
        7618 => x"00000016", -- pedding 
        7619 => x"00000016", -- pedding 
        7620 => x"00000016", -- pedding 
        7621 => x"00000016", -- pedding 
        7622 => x"00000016", -- pedding 
        7623 => x"00000016", -- pedding 
        7624 => x"00000016", -- pedding 
        7625 => x"00000016", -- pedding 
        7626 => x"00000016", -- pedding 
        7627 => x"00000016", -- pedding 
        7628 => x"00000016", -- pedding 
        7629 => x"00000016", -- pedding 
        7630 => x"00000016", -- pedding 
        7631 => x"00000016", -- pedding 
        7632 => x"00000016", -- pedding 
        7633 => x"00000016", -- pedding 
        7634 => x"00000016", -- pedding 
        7635 => x"00000016", -- pedding 
        7636 => x"00000016", -- pedding 
        7637 => x"00000016", -- pedding 
        7638 => x"00000016", -- pedding 
        7639 => x"00000016", -- pedding 
        7640 => x"00000016", -- pedding 
        7641 => x"00000016", -- pedding 
        7642 => x"00000016", -- pedding 
        7643 => x"00000016", -- pedding 
        7644 => x"00000016", -- pedding 
        7645 => x"00000016", -- pedding 
        7646 => x"00000016", -- pedding 
        7647 => x"00000016", -- pedding 
        7648 => x"00000016", -- pedding 
        7649 => x"00000016", -- pedding 
        7650 => x"00000016", -- pedding 
        7651 => x"00000016", -- pedding 
        7652 => x"00000016", -- pedding 
        7653 => x"00000016", -- pedding 
        7654 => x"00000016", -- pedding 
        7655 => x"00000016", -- pedding 
        7656 => x"00000016", -- pedding 
        7657 => x"00000016", -- pedding 
        7658 => x"00000016", -- pedding 
        7659 => x"00000016", -- pedding 
        7660 => x"00000016", -- pedding 
        7661 => x"00000016", -- pedding 
        7662 => x"00000016", -- pedding 
        7663 => x"00000016", -- pedding 
        7664 => x"00000016", -- pedding 
        7665 => x"00000016", -- pedding 
        7666 => x"00000016", -- pedding 
        7667 => x"00000016", -- pedding 
        7668 => x"00000016", -- pedding 
        7669 => x"00000016", -- pedding 
        7670 => x"00000016", -- pedding 
        7671 => x"00000016", -- pedding 
        7672 => x"00000016", -- pedding 
        7673 => x"00000016", -- pedding 
        7674 => x"00000016", -- pedding 
        7675 => x"00000016", -- pedding 
        7676 => x"00000016", -- pedding 
        7677 => x"00000016", -- pedding 
        7678 => x"00000016", -- pedding 
        7679 => x"00000016", -- pedding 
        7680 => x"00000016", -- pedding 
        7681 => x"00000016", -- pedding 
        7682 => x"00000016", -- pedding 
        7683 => x"00000016", -- pedding 
        7684 => x"00000016", -- pedding 
        7685 => x"00000016", -- pedding 
        7686 => x"00000016", -- pedding 
        7687 => x"00000016", -- pedding 
        7688 => x"00000016", -- pedding 
        7689 => x"00000016", -- pedding 
        7690 => x"00000016", -- pedding 
        7691 => x"00000016", -- pedding 
        7692 => x"00000016", -- pedding 
        7693 => x"00000016", -- pedding 
        7694 => x"00000016", -- pedding 
        7695 => x"00000016", -- pedding 
        7696 => x"00000016", -- pedding 
        7697 => x"00000016", -- pedding 
        7698 => x"00000016", -- pedding 
        7699 => x"00000016", -- pedding 
        7700 => x"00000016", -- pedding 
        7701 => x"00000016", -- pedding 
        7702 => x"00000016", -- pedding 
        7703 => x"00000016", -- pedding 
        7704 => x"00000016", -- pedding 
        7705 => x"00000016", -- pedding 
        7706 => x"00000016", -- pedding 
        7707 => x"00000016", -- pedding 
        7708 => x"00000016", -- pedding 
        7709 => x"00000016", -- pedding 
        7710 => x"00000016", -- pedding 
        7711 => x"00000016", -- pedding 
        7712 => x"00000016", -- pedding 
        7713 => x"00000016", -- pedding 
        7714 => x"00000016", -- pedding 
        7715 => x"00000016", -- pedding 
        7716 => x"00000016", -- pedding 
        7717 => x"00000016", -- pedding 
        7718 => x"00000016", -- pedding 
        7719 => x"00000016", -- pedding 
        7720 => x"00000016", -- pedding 
        7721 => x"00000016", -- pedding 
        7722 => x"00000016", -- pedding 
        7723 => x"00000016", -- pedding 
        7724 => x"00000016", -- pedding 
        7725 => x"00000016", -- pedding 
        7726 => x"00000016", -- pedding 
        7727 => x"00000016", -- pedding 
        7728 => x"00000016", -- pedding 
        7729 => x"00000016", -- pedding 
        7730 => x"00000016", -- pedding 
        7731 => x"00000016", -- pedding 
        7732 => x"00000016", -- pedding 
        7733 => x"00000016", -- pedding 
        7734 => x"00000016", -- pedding 
        7735 => x"00000016", -- pedding 
        7736 => x"00000016", -- pedding 
        7737 => x"00000016", -- pedding 
        7738 => x"00000016", -- pedding 
        7739 => x"00000016", -- pedding 
        7740 => x"00000016", -- pedding 
        7741 => x"00000016", -- pedding 
        7742 => x"00000016", -- pedding 
        7743 => x"00000016", -- pedding 
        7744 => x"00000016", -- pedding 
        7745 => x"00000016", -- pedding 
        7746 => x"00000016", -- pedding 
        7747 => x"00000016", -- pedding 
        7748 => x"00000016", -- pedding 
        7749 => x"00000016", -- pedding 
        7750 => x"00000016", -- pedding 
        7751 => x"00000016", -- pedding 
        7752 => x"00000016", -- pedding 
        7753 => x"00000016", -- pedding 
        7754 => x"00000016", -- pedding 
        7755 => x"00000016", -- pedding 
        7756 => x"00000016", -- pedding 
        7757 => x"00000016", -- pedding 
        7758 => x"00000016", -- pedding 
        7759 => x"00000016", -- pedding 
        7760 => x"00000016", -- pedding 
        7761 => x"00000016", -- pedding 
        7762 => x"00000016", -- pedding 
        7763 => x"00000016", -- pedding 
        7764 => x"00000016", -- pedding 
        7765 => x"00000016", -- pedding 
        7766 => x"00000016", -- pedding 
        7767 => x"00000016", -- pedding 
        7768 => x"00000016", -- pedding 
        7769 => x"00000016", -- pedding 
        7770 => x"00000016", -- pedding 
        7771 => x"00000016", -- pedding 
        7772 => x"00000016", -- pedding 
        7773 => x"00000016", -- pedding 
        7774 => x"00000016", -- pedding 
        7775 => x"00000016", -- pedding 
        7776 => x"00000016", -- pedding 
        7777 => x"00000016", -- pedding 
        7778 => x"00000016", -- pedding 
        7779 => x"00000016", -- pedding 
        7780 => x"00000016", -- pedding 
        7781 => x"00000016", -- pedding 
        7782 => x"00000016", -- pedding 
        7783 => x"00000016", -- pedding 
        7784 => x"00000016", -- pedding 
        7785 => x"00000016", -- pedding 
        7786 => x"00000016", -- pedding 
        7787 => x"00000016", -- pedding 
        7788 => x"00000016", -- pedding 
        7789 => x"00000016", -- pedding 
        7790 => x"00000016", -- pedding 
        7791 => x"00000016", -- pedding 
        7792 => x"00000016", -- pedding 
        7793 => x"00000016", -- pedding 
        7794 => x"00000016", -- pedding 
        7795 => x"00000016", -- pedding 
        7796 => x"00000016", -- pedding 
        7797 => x"00000016", -- pedding 
        7798 => x"00000016", -- pedding 
        7799 => x"00000016", -- pedding 
        7800 => x"00000016", -- pedding 
        7801 => x"00000016", -- pedding 
        7802 => x"00000016", -- pedding 
        7803 => x"00000016", -- pedding 
        7804 => x"00000016", -- pedding 
        7805 => x"00000016", -- pedding 
        7806 => x"00000016", -- pedding 
        7807 => x"00000016", -- pedding 
        7808 => x"00000016", -- pedding 
        7809 => x"00000016", -- pedding 
        7810 => x"00000016", -- pedding 
        7811 => x"00000016", -- pedding 
        7812 => x"00000016", -- pedding 
        7813 => x"00000016", -- pedding 
        7814 => x"00000016", -- pedding 
        7815 => x"00000016", -- pedding 
        7816 => x"00000016", -- pedding 
        7817 => x"00000016", -- pedding 
        7818 => x"00000016", -- pedding 
        7819 => x"00000016", -- pedding 
        7820 => x"00000016", -- pedding 
        7821 => x"00000016", -- pedding 
        7822 => x"00000016", -- pedding 
        7823 => x"00000016", -- pedding 
        7824 => x"00000016", -- pedding 
        7825 => x"00000016", -- pedding 
        7826 => x"00000016", -- pedding 
        7827 => x"00000016", -- pedding 
        7828 => x"00000016", -- pedding 
        7829 => x"00000016", -- pedding 
        7830 => x"00000016", -- pedding 
        7831 => x"00000016", -- pedding 
        7832 => x"00000016", -- pedding 
        7833 => x"00000016", -- pedding 
        7834 => x"00000016", -- pedding 
        7835 => x"00000016", -- pedding 
        7836 => x"00000016", -- pedding 
        7837 => x"00000016", -- pedding 
        7838 => x"00000016", -- pedding 
        7839 => x"00000016", -- pedding 
        7840 => x"00000016", -- pedding 
        7841 => x"00000016", -- pedding 
        7842 => x"00000016", -- pedding 
        7843 => x"00000016", -- pedding 
        7844 => x"00000016", -- pedding 
        7845 => x"00000016", -- pedding 
        7846 => x"00000016", -- pedding 
        7847 => x"00000016", -- pedding 
        7848 => x"00000016", -- pedding 
        7849 => x"00000016", -- pedding 
        7850 => x"00000016", -- pedding 
        7851 => x"00000016", -- pedding 
        7852 => x"00000016", -- pedding 
        7853 => x"00000016", -- pedding 
        7854 => x"00000016", -- pedding 
        7855 => x"00000016", -- pedding 
        7856 => x"00000016", -- pedding 
        7857 => x"00000016", -- pedding 
        7858 => x"00000016", -- pedding 
        7859 => x"00000016", -- pedding 
        7860 => x"00000016", -- pedding 
        7861 => x"00000016", -- pedding 
        7862 => x"00000016", -- pedding 
        7863 => x"00000016", -- pedding 
        7864 => x"00000016", -- pedding 
        7865 => x"00000016", -- pedding 
        7866 => x"00000016", -- pedding 
        7867 => x"00000016", -- pedding 
        7868 => x"00000016", -- pedding 
        7869 => x"00000016", -- pedding 
        7870 => x"00000016", -- pedding 
        7871 => x"00000016", -- pedding 
        7872 => x"00000016", -- pedding 
        7873 => x"00000016", -- pedding 
        7874 => x"00000016", -- pedding 
        7875 => x"00000016", -- pedding 
        7876 => x"00000016", -- pedding 
        7877 => x"00000016", -- pedding 
        7878 => x"00000016", -- pedding 
        7879 => x"00000016", -- pedding 
        7880 => x"00000016", -- pedding 
        7881 => x"00000016", -- pedding 
        7882 => x"00000016", -- pedding 
        7883 => x"00000016", -- pedding 
        7884 => x"00000016", -- pedding 
        7885 => x"00000016", -- pedding 
        7886 => x"00000016", -- pedding 
        7887 => x"00000016", -- pedding 
        7888 => x"00000016", -- pedding 
        7889 => x"00000016", -- pedding 
        7890 => x"00000016", -- pedding 
        7891 => x"00000016", -- pedding 
        7892 => x"00000016", -- pedding 
        7893 => x"00000016", -- pedding 
        7894 => x"00000016", -- pedding 
        7895 => x"00000016", -- pedding 
        7896 => x"00000016", -- pedding 
        7897 => x"00000016", -- pedding 
        7898 => x"00000016", -- pedding 
        7899 => x"00000016", -- pedding 
        7900 => x"00000016", -- pedding 
        7901 => x"00000016", -- pedding 
        7902 => x"00000016", -- pedding 
        7903 => x"00000016", -- pedding 
        7904 => x"00000016", -- pedding 
        7905 => x"00000016", -- pedding 
        7906 => x"00000016", -- pedding 
        7907 => x"00000016", -- pedding 
        7908 => x"00000016", -- pedding 
        7909 => x"00000016", -- pedding 
        7910 => x"00000016", -- pedding 
        7911 => x"00000016", -- pedding 
        7912 => x"00000016", -- pedding 
        7913 => x"00000016", -- pedding 
        7914 => x"00000016", -- pedding 
        7915 => x"00000016", -- pedding 
        7916 => x"00000016", -- pedding 
        7917 => x"00000016", -- pedding 
        7918 => x"00000016", -- pedding 
        7919 => x"00000016", -- pedding 
        7920 => x"00000016", -- pedding 
        7921 => x"00000016", -- pedding 
        7922 => x"00000016", -- pedding 
        7923 => x"00000016", -- pedding 
        7924 => x"00000016", -- pedding 
        7925 => x"00000016", -- pedding 
        7926 => x"00000016", -- pedding 
        7927 => x"00000016", -- pedding 
        7928 => x"00000016", -- pedding 
        7929 => x"00000016", -- pedding 
        7930 => x"00000016", -- pedding 
        7931 => x"00000016", -- pedding 
        7932 => x"00000016", -- pedding 
        7933 => x"00000016", -- pedding 
        7934 => x"00000016", -- pedding 
        7935 => x"00000016", -- pedding 
        7936 => x"00000016", -- pedding 
        7937 => x"00000016", -- pedding 
        7938 => x"00000016", -- pedding 
        7939 => x"00000016", -- pedding 
        7940 => x"00000016", -- pedding 
        7941 => x"00000016", -- pedding 
        7942 => x"00000016", -- pedding 
        7943 => x"00000016", -- pedding 
        7944 => x"00000016", -- pedding 
        7945 => x"00000016", -- pedding 
        7946 => x"00000016", -- pedding 
        7947 => x"00000016", -- pedding 
        7948 => x"00000016", -- pedding 
        7949 => x"00000016", -- pedding 
        7950 => x"00000016", -- pedding 
        7951 => x"00000016", -- pedding 
        7952 => x"00000016", -- pedding 
        7953 => x"00000016", -- pedding 
        7954 => x"00000016", -- pedding 
        7955 => x"00000016", -- pedding 
        7956 => x"00000016", -- pedding 
        7957 => x"00000016", -- pedding 
        7958 => x"00000016", -- pedding 
        7959 => x"00000016", -- pedding 
        7960 => x"00000016", -- pedding 
        7961 => x"00000016", -- pedding 
        7962 => x"00000016", -- pedding 
        7963 => x"00000016", -- pedding 
        7964 => x"00000016", -- pedding 
        7965 => x"00000016", -- pedding 
        7966 => x"00000016", -- pedding 
        7967 => x"00000016", -- pedding 
        7968 => x"00000016", -- pedding 
        7969 => x"00000016", -- pedding 
        7970 => x"00000016", -- pedding 
        7971 => x"00000016", -- pedding 
        7972 => x"00000016", -- pedding 
        7973 => x"00000016", -- pedding 
        7974 => x"00000016", -- pedding 
        7975 => x"00000016", -- pedding 
        7976 => x"00000016", -- pedding 
        7977 => x"00000016", -- pedding 
        7978 => x"00000016", -- pedding 
        7979 => x"00000016", -- pedding 
        7980 => x"00000016", -- pedding 
        7981 => x"00000016", -- pedding 
        7982 => x"00000016", -- pedding 
        7983 => x"00000016", -- pedding 
        7984 => x"00000016", -- pedding 
        7985 => x"00000016", -- pedding 
        7986 => x"00000016", -- pedding 
        7987 => x"00000016", -- pedding 
        7988 => x"00000016", -- pedding 
        7989 => x"00000016", -- pedding 
        7990 => x"00000016", -- pedding 
        7991 => x"00000016", -- pedding 
        7992 => x"00000016", -- pedding 
        7993 => x"00000016", -- pedding 
        7994 => x"00000016", -- pedding 
        7995 => x"00000016", -- pedding 
        7996 => x"00000016", -- pedding 
        7997 => x"00000016", -- pedding 
        7998 => x"00000016", -- pedding 
        7999 => x"00000016", -- pedding 
        8000 => x"00000016", -- pedding 
        8001 => x"00000016", -- pedding 
        8002 => x"00000016", -- pedding 
        8003 => x"00000016", -- pedding 
        8004 => x"00000016", -- pedding 
        8005 => x"00000016", -- pedding 
        8006 => x"00000016", -- pedding 
        8007 => x"00000016", -- pedding 
        8008 => x"00000016", -- pedding 
        8009 => x"00000016", -- pedding 
        8010 => x"00000016", -- pedding 
        8011 => x"00000016", -- pedding 
        8012 => x"00000016", -- pedding 
        8013 => x"00000016", -- pedding 
        8014 => x"00000016", -- pedding 
        8015 => x"00000016", -- pedding 
        8016 => x"00000016", -- pedding 
        8017 => x"00000016", -- pedding 
        8018 => x"00000016", -- pedding 
        8019 => x"00000016", -- pedding 
        8020 => x"00000016", -- pedding 
        8021 => x"00000016", -- pedding 
        8022 => x"00000016", -- pedding 
        8023 => x"00000016", -- pedding 
        8024 => x"00000016", -- pedding 
        8025 => x"00000016", -- pedding 
        8026 => x"00000016", -- pedding 
        8027 => x"00000016", -- pedding 
        8028 => x"00000016", -- pedding 
        8029 => x"00000016", -- pedding 
        8030 => x"00000016", -- pedding 
        8031 => x"00000016", -- pedding 
        8032 => x"00000016", -- pedding 
        8033 => x"00000016", -- pedding 
        8034 => x"00000016", -- pedding 
        8035 => x"00000016", -- pedding 
        8036 => x"00000016", -- pedding 
        8037 => x"00000016", -- pedding 
        8038 => x"00000016", -- pedding 
        8039 => x"00000016", -- pedding 
        8040 => x"00000016", -- pedding 
        8041 => x"00000016", -- pedding 
        8042 => x"00000016", -- pedding 
        8043 => x"00000016", -- pedding 
        8044 => x"00000016", -- pedding 
        8045 => x"00000016", -- pedding 
        8046 => x"00000016", -- pedding 
        8047 => x"00000016", -- pedding 
        8048 => x"00000016", -- pedding 
        8049 => x"00000016", -- pedding 
        8050 => x"00000016", -- pedding 
        8051 => x"00000016", -- pedding 
        8052 => x"00000016", -- pedding 
        8053 => x"00000016", -- pedding 
        8054 => x"00000016", -- pedding 
        8055 => x"00000016", -- pedding 
        8056 => x"00000016", -- pedding 
        8057 => x"00000016", -- pedding 
        8058 => x"00000016", -- pedding 
        8059 => x"00000016", -- pedding 
        8060 => x"00000016", -- pedding 
        8061 => x"00000016", -- pedding 
        8062 => x"00000016", -- pedding 
        8063 => x"00000016", -- pedding 
        8064 => x"00000016", -- pedding 
        8065 => x"00000016", -- pedding 
        8066 => x"00000016", -- pedding 
        8067 => x"00000016", -- pedding 
        8068 => x"00000016", -- pedding 
        8069 => x"00000016", -- pedding 
        8070 => x"00000016", -- pedding 
        8071 => x"00000016", -- pedding 
        8072 => x"00000016", -- pedding 
        8073 => x"00000016", -- pedding 
        8074 => x"00000016", -- pedding 
        8075 => x"00000016", -- pedding 
        8076 => x"00000016", -- pedding 
        8077 => x"00000016", -- pedding 
        8078 => x"00000016", -- pedding 
        8079 => x"00000016", -- pedding 
        8080 => x"00000016", -- pedding 
        8081 => x"00000016", -- pedding 
        8082 => x"00000016", -- pedding 
        8083 => x"00000016", -- pedding 
        8084 => x"00000016", -- pedding 
        8085 => x"00000016", -- pedding 
        8086 => x"00000016", -- pedding 
        8087 => x"00000016", -- pedding 
        8088 => x"00000016", -- pedding 
        8089 => x"00000016", -- pedding 
        8090 => x"00000016", -- pedding 
        8091 => x"00000016", -- pedding 
        8092 => x"00000016", -- pedding 
        8093 => x"00000016", -- pedding 
        8094 => x"00000016", -- pedding 
        8095 => x"00000016", -- pedding 
        8096 => x"00000016", -- pedding 
        8097 => x"00000016", -- pedding 
        8098 => x"00000016", -- pedding 
        8099 => x"00000016", -- pedding 
others => x"00000000"
	);


begin

	process(i_clk)
	begin
		if rising_edge(i_clk) then
			-- memory write --
			if i_we = '1' then
				mem(to_integer(unsigned(i_w_addr))) <= i_data;
			end if;
			-- memory read -- 
			o_data <= mem(to_integer(unsigned(i_r_addr)));
			
		end if; 
	end process;

end architecture arch;
