
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity ram is
	generic
	(
		DATA_WIDTH : natural := 32;		    -- 4 byte one line of memory
		ADDR_WIDTH : natural := 13			    -- 24576 bytes size of memory
	);

	port(
		i_clk    : in  std_logic;
		i_r_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		i_data   : in  std_logic_vector(DATA_WIDTH-1 downto 0);
		i_we     : in  std_logic;
		i_w_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		o_data   : out std_logic_vector(DATA_WIDTH-1 downto 0)
	);
end entity ram;

architecture arch of ram is

	type ram_t is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(DATA_WIDTH-1 downto 0);


-- GENERATED BY BC_MEM_PACKER

-- DATE: Thu May 18 16:01:02 2017

	signal mem : ram_t := (

--			***** COLOR PALLETE *****

		-- fellas
		0 =>	x"00C84C0C", -- R: 0 G: 0 B: 0
		1 =>	x"00FCD8A8", -- R: 222 G: 89 B: 24
		2 =>	x"00000000", -- R: 255 G: 242 B: 226
		3 =>	x"002038EC", -- R: 0 G: 162 B: 232
		4 =>	x"0000A800", -- R: 251 G: 157 B: 66
		5 =>	x"00FCFCFC", -- R: 252 G: 150 B: 52
		6 =>	x"00747474", -- R: 255 G: 157 B: 58
		7 =>	x"00C0C0C0", -- R: 255 G: 157 B: 59
		--below not fellas
		8 =>	x"003599FF", -- R: 255 G: 153 B: 53
		9 =>	x"004B91C0", -- R: 192 G: 145 B: 75
		10 =>	x"00947C00", -- R: 0 G: 124 B: 148
		11 =>	x"00877D00", -- R: 0 G: 125 B: 135
		12 =>	x"008E860E", -- R: 14 G: 134 B: 142
		13 =>	x"003B9AFC", -- R: 252 G: 154 B: 59
		14 =>	x"00399DFF", -- R: 255 G: 157 B: 57
		15 =>	x"001C68DB", -- R: 219 G: 104 B: 28
		16 =>	x"001E6CDE", -- R: 222 G: 108 B: 30
		17 =>	x"003495FF", -- R: 255 G: 149 B: 52
		18 =>	x"003F96E6", -- R: 230 G: 150 B: 63
		19 =>	x"005A8D8E", -- R: 142 G: 141 B: 90
		20 =>	x"007C821E", -- R: 30 G: 130 B: 124
		21 =>	x"008C8100", -- R: 0 G: 129 B: 140
		22 =>	x"00208BFB", -- R: 251 G: 139 B: 32
		23 =>	x"003697FC", -- R: 252 G: 151 B: 54
		24 =>	x"003CA0FF", -- R: 255 G: 160 B: 60
		25 =>	x"000540C0", -- R: 192 G: 64 B: 5
		26 =>	x"000846C4", -- R: 196 G: 70 B: 8
		27 =>	x"00043FC1", -- R: 193 G: 63 B: 4
		28 =>	x"003491F7", -- R: 247 G: 145 B: 52
		29 =>	x"003799FF", -- R: 255 G: 153 B: 55
		30 =>	x"002C9BFF", -- R: 255 G: 155 B: 44
		31 =>	x"00728640", -- R: 64 G: 134 B: 114
		32 =>	x"00897E00", -- R: 0 G: 126 B: 137
		33 =>	x"007A7000", -- R: 0 G: 112 B: 122
		34 =>	x"00218CFB", -- R: 251 G: 140 B: 33
		35 =>	x"002B91FB", -- R: 251 G: 145 B: 43
		36 =>	x"001C68DA", -- R: 218 G: 104 B: 28
		37 =>	x"000035B8", -- R: 184 G: 53 B: 0
		38 =>	x"0041A8FF", -- R: 255 G: 168 B: 65
		39 =>	x"003DA0FF", -- R: 255 G: 160 B: 61
		40 =>	x"0034A3FF", -- R: 255 G: 163 B: 52
		41 =>	x"008C8000", -- R: 0 G: 128 B: 140
		42 =>	x"007E831C", -- R: 28 G: 131 B: 126
		43 =>	x"00309AFF", -- R: 255 G: 154 B: 48
		44 =>	x"003399FF", -- R: 255 G: 153 B: 51
		45 =>	x"00577AB9", -- R: 185 G: 122 B: 87
		46 =>	x"00807700", -- R: 0 G: 119 B: 128
		47 =>	x"007A7100", -- R: 0 G: 113 B: 122
		48 =>	x"003898FC", -- R: 252 G: 152 B: 56
		49 =>	x"001F6DDE", -- R: 222 G: 109 B: 31
		50 =>	x"00043EBE", -- R: 190 G: 62 B: 4
		51 =>	x"002F9AFF", -- R: 255 G: 154 B: 47
		52 =>	x"00848109", -- R: 9 G: 129 B: 132
		53 =>	x"003698FF", -- R: 255 G: 152 B: 54
		54 =>	x"003B97EF", -- R: 239 G: 151 B: 59
		55 =>	x"0033A2FF", -- R: 255 G: 162 B: 51
		56 =>	x"00269DFF", -- R: 255 G: 157 B: 38
		57 =>	x"008A7F00", -- R: 0 G: 127 B: 138
		58 =>	x"002E9AFF", -- R: 255 G: 154 B: 46
		59 =>	x"008D7E00", -- R: 0 G: 126 B: 141
		60 =>	x"003F95E4", -- R: 228 G: 149 B: 63
		61 =>	x"003598FF", -- R: 255 G: 152 B: 53
		62 =>	x"003C9AFC", -- R: 252 G: 154 B: 60
		63 =>	x"003199FF", -- R: 255 G: 153 B: 49
		64 =>	x"0069885F", -- R: 95 G: 136 B: 105
		65 =>	x"00658A6C", -- R: 108 G: 138 B: 101
		66 =>	x"006A895E", -- R: 94 G: 137 B: 106
		67 =>	x"003997F7", -- R: 247 G: 151 B: 57
		68 =>	x"003E95E8", -- R: 232 G: 149 B: 62
		69 =>	x"003299FF", -- R: 255 G: 153 B: 50
		70 =>	x"003499FF", -- R: 255 G: 153 B: 52
		71 =>	x"004A91C0", -- R: 192 G: 145 B: 74
		72 =>	x"00277FFF", -- R: 255 G: 127 B: 39
		73 =>	x"00584000", -- R: 0 G: 64 B: 88
		74 =>	x"00C9DDFF", -- R: 255 G: 221 B: 201
		75 =>	x"000038F8", -- R: 248 G: 56 B: 0
		76 =>	x"00007CAC", -- R: 172 G: 124 B: 0
		77 =>	x"0040A4FF", -- R: 255 G: 164 B: 64
		78 =>	x"00349DEF", -- R: 239 G: 157 B: 52
		79 =>	x"003092E0", -- R: 224 G: 146 B: 48
		80 =>	x"00309AEA", -- R: 234 G: 154 B: 48
		81 =>	x"00000000", -- Unused
		82 =>	x"00000000", -- Unused
		83 =>	x"00000000", -- Unused
		84 =>	x"00000000", -- Unused
		85 =>	x"00000000", -- Unused
		86 =>	x"00000000", -- Unused
		87 =>	x"00000000", -- Unused
		88 =>	x"00000000", -- Unused
		89 =>	x"00000000", -- Unused
		90 =>	x"00000000", -- Unused
		91 =>	x"00000000", -- Unused
		92 =>	x"00000000", -- Unused
		93 =>	x"00000000", -- Unused
		94 =>	x"00000000", -- Unused
		95 =>	x"00000000", -- Unused
		96 =>	x"00000000", -- Unused
		97 =>	x"00000000", -- Unused
		98 =>	x"00000000", -- Unused
		99 =>	x"00000000", -- Unused
		100 =>	x"00000000", -- Unused
		101 =>	x"00000000", -- Unused
		102 =>	x"00000000", -- Unused
		103 =>	x"00000000", -- Unused
		104 =>	x"00000000", -- Unused
		105 =>	x"00000000", -- Unused
		106 =>	x"00000000", -- Unused
		107 =>	x"00000000", -- Unused
		108 =>	x"00000000", -- Unused
		109 =>	x"00000000", -- Unused
		110 =>	x"00000000", -- Unused
		111 =>	x"00000000", -- Unused
		112 =>	x"00000000", -- Unused
		113 =>	x"00000000", -- Unused
		114 =>	x"00000000", -- Unused
		115 =>	x"00000000", -- Unused
		116 =>	x"00000000", -- Unused
		117 =>	x"00000000", -- Unused
		118 =>	x"00000000", -- Unused
		119 =>	x"00000000", -- Unused
		120 =>	x"00000000", -- Unused
		121 =>	x"00000000", -- Unused
		122 =>	x"00000000", -- Unused
		123 =>	x"00000000", -- Unused
		124 =>	x"00000000", -- Unused
		125 =>	x"00000000", -- Unused
		126 =>	x"00000000", -- Unused
		127 =>	x"00000000", -- Unused
		128 =>	x"00000000", -- Unused
		129 =>	x"00000000", -- Unused
		130 =>	x"00000000", -- Unused
		131 =>	x"00000000", -- Unused
		132 =>	x"00000000", -- Unused
		133 =>	x"00000000", -- Unused
		134 =>	x"00000000", -- Unused
		135 =>	x"00000000", -- Unused
		136 =>	x"00000000", -- Unused
		137 =>	x"00000000", -- Unused
		138 =>	x"00000000", -- Unused
		139 =>	x"00000000", -- Unused
		140 =>	x"00000000", -- Unused
		141 =>	x"00000000", -- Unused
		142 =>	x"00000000", -- Unused
		143 =>	x"00000000", -- Unused
		144 =>	x"00000000", -- Unused
		145 =>	x"00000000", -- Unused
		146 =>	x"00000000", -- Unused
		147 =>	x"00000000", -- Unused
		148 =>	x"00000000", -- Unused
		149 =>	x"00000000", -- Unused
		150 =>	x"00000000", -- Unused
		151 =>	x"00000000", -- Unused
		152 =>	x"00000000", -- Unused
		153 =>	x"00000000", -- Unused
		154 =>	x"00000000", -- Unused
		155 =>	x"00000000", -- Unused
		156 =>	x"00000000", -- Unused
		157 =>	x"00000000", -- Unused
		158 =>	x"00000000", -- Unused
		159 =>	x"00000000", -- Unused
		160 =>	x"00000000", -- Unused
		161 =>	x"00000000", -- Unused
		162 =>	x"00000000", -- Unused
		163 =>	x"00000000", -- Unused
		164 =>	x"00000000", -- Unused
		165 =>	x"00000000", -- Unused
		166 =>	x"00000000", -- Unused
		167 =>	x"00000000", -- Unused
		168 =>	x"00000000", -- Unused
		169 =>	x"00000000", -- Unused
		170 =>	x"00000000", -- Unused
		171 =>	x"00000000", -- Unused
		172 =>	x"00000000", -- Unused
		173 =>	x"00000000", -- Unused
		174 =>	x"00000000", -- Unused
		175 =>	x"00000000", -- Unused
		176 =>	x"00000000", -- Unused
		177 =>	x"00000000", -- Unused
		178 =>	x"00000000", -- Unused
		179 =>	x"00000000", -- Unused
		180 =>	x"00000000", -- Unused
		181 =>	x"00000000", -- Unused
		182 =>	x"00000000", -- Unused
		183 =>	x"00000000", -- Unused
		184 =>	x"00000000", -- Unused
		185 =>	x"00000000", -- Unused
		186 =>	x"00000000", -- Unused
		187 =>	x"00000000", -- Unused
		188 =>	x"00000000", -- Unused
		189 =>	x"00000000", -- Unused
		190 =>	x"00000000", -- Unused
		191 =>	x"00000000", -- Unused
		192 =>	x"00000000", -- Unused
		193 =>	x"00000000", -- Unused
		194 =>	x"00000000", -- Unused
		195 =>	x"00000000", -- Unused
		196 =>	x"00000000", -- Unused
		197 =>	x"00000000", -- Unused
		198 =>	x"00000000", -- Unused
		199 =>	x"00000000", -- Unused
		200 =>	x"00000000", -- Unused
		201 =>	x"00000000", -- Unused
		202 =>	x"00000000", -- Unused
		203 =>	x"00000000", -- Unused
		204 =>	x"00000000", -- Unused
		205 =>	x"00000000", -- Unused
		206 =>	x"00000000", -- Unused
		207 =>	x"00000000", -- Unused
		208 =>	x"00000000", -- Unused
		209 =>	x"00000000", -- Unused
		210 =>	x"00000000", -- Unused
		211 =>	x"00000000", -- Unused
		212 =>	x"00000000", -- Unused
		213 =>	x"00000000", -- Unused
		214 =>	x"00000000", -- Unused
		215 =>	x"00000000", -- Unused
		216 =>	x"00000000", -- Unused
		217 =>	x"00000000", -- Unused
		218 =>	x"00000000", -- Unused
		219 =>	x"00000000", -- Unused
		220 =>	x"00000000", -- Unused
		221 =>	x"00000000", -- Unused
		222 =>	x"00000000", -- Unused
		223 =>	x"00000000", -- Unused
		224 =>	x"00000000", -- Unused
		225 =>	x"00000000", -- Unused
		226 =>	x"00000000", -- Unused
		227 =>	x"00000000", -- Unused
		228 =>	x"00000000", -- Unused
		229 =>	x"00000000", -- Unused
		230 =>	x"00000000", -- Unused
		231 =>	x"00000000", -- Unused
		232 =>	x"00000000", -- Unused
		233 =>	x"00000000", -- Unused
		234 =>	x"00000000", -- Unused
		235 =>	x"00000000", -- Unused
		236 =>	x"00000000", -- Unused
		237 =>	x"00000000", -- Unused
		238 =>	x"00000000", -- Unused
		239 =>	x"00000000", -- Unused
		240 =>	x"00000000", -- Unused
		241 =>	x"00000000", -- Unused
		242 =>	x"00000000", -- Unused
		243 =>	x"00000000", -- Unused
		244 =>	x"00000000", -- Unused
		245 =>	x"00000000", -- Unused
		246 =>	x"00000000", -- Unused
		247 =>	x"00000000", -- Unused
		248 =>	x"00000000", -- Unused
		249 =>	x"00000000", -- Unused
		250 =>	x"00000000", -- Unused
		251 =>	x"00000000", -- Unused
		252 =>	x"00000000", -- Unused
		253 =>	x"00000000", -- Unused
		254 =>	x"00000000", -- Unused

--			***** 16x16 IMAGES *****
                --  sprite 0
        255 => x"00000000",
        256 => x"00000000",
        257 => x"00000000",
        258 => x"00000000",
        259 => x"01010000",
        260 => x"02010101",
        261 => x"01010101",
        262 => x"01010101",
        263 => x"01010101",
        264 => x"01010101",
        265 => x"01010101",
        266 => x"01010101",
        267 => x"01000101",
        268 => x"01030301",
        269 => x"01010100",
        270 => x"01010101",
        271 => x"01020202",
        272 => x"02010101",
        273 => x"01020202",
        274 => x"02020201",
        275 => x"01010101",
        276 => x"01010201",
        277 => x"01010101",
        278 => x"01010101",
        279 => x"04040404",
        280 => x"04040404",
        281 => x"04040404",
        282 => x"04040404",
        283 => x"01010404",
        284 => x"02010101",
        285 => x"01010101",
        286 => x"01010101",
        287 => x"01010101",
        288 => x"01010101",
        289 => x"01010101",
        290 => x"01010101",
        291 => x"01040101",
        292 => x"01030301",
        293 => x"01010104",
        294 => x"01010101",
        295 => x"01020202",
        296 => x"02010101",
        297 => x"01020202",
        298 => x"02020201",
        299 => x"01010101",
        300 => x"01010201",
        301 => x"01010101",
        302 => x"01010101",
        303 => x"05050505",
        304 => x"05050505",
        305 => x"05050505",
        306 => x"05050505",
        307 => x"06060505",
        308 => x"02060606",
        309 => x"06060606",
        310 => x"06060606",
        311 => x"06060606",
        312 => x"06060606",
        313 => x"06060606",
        314 => x"06060606",
        315 => x"06050606",
        316 => x"06030306",
        317 => x"06060605",
        318 => x"06060606",
        319 => x"06020202",
        320 => x"02060606",
        321 => x"06020202",
        322 => x"02020206",
        323 => x"06060606",
        324 => x"06060206",
        325 => x"06060606",
        326 => x"06060606",

                --  sprite 1
        327 => x"00020202",
        328 => x"02020202",
        329 => x"02020202",
        330 => x"02020200",
        331 => x"01000000",
        332 => x"00020101",
        333 => x"01010101",
        334 => x"01010101",
        335 => x"01010101",
        336 => x"01010101",
        337 => x"01010101",
        338 => x"01010101",
        339 => x"01000000",
        340 => x"03030303",
        341 => x"01010100",
        342 => x"00020202",
        343 => x"02020202",
        344 => x"02020101",
        345 => x"02020202",
        346 => x"02020202",
        347 => x"01010101",
        348 => x"01020201",
        349 => x"01010101",
        350 => x"01010101",
        351 => x"04020202",
        352 => x"02020202",
        353 => x"02020202",
        354 => x"02020204",
        355 => x"01040404",
        356 => x"04020101",
        357 => x"01010101",
        358 => x"01010101",
        359 => x"01010101",
        360 => x"01010101",
        361 => x"01010101",
        362 => x"01010101",
        363 => x"01040404",
        364 => x"03030303",
        365 => x"01010104",
        366 => x"04020202",
        367 => x"02020202",
        368 => x"02020101",
        369 => x"02020202",
        370 => x"02020202",
        371 => x"01010101",
        372 => x"01020201",
        373 => x"01010101",
        374 => x"01010101",
        375 => x"05020202",
        376 => x"02020202",
        377 => x"02020202",
        378 => x"02020205",
        379 => x"06050505",
        380 => x"05020606",
        381 => x"06060606",
        382 => x"06060606",
        383 => x"06060606",
        384 => x"06060606",
        385 => x"06060606",
        386 => x"06060606",
        387 => x"06050505",
        388 => x"03030303",
        389 => x"06060605",
        390 => x"05020202",
        391 => x"02020202",
        392 => x"02020606",
        393 => x"02020202",
        394 => x"02020202",
        395 => x"06060606",
        396 => x"06020206",
        397 => x"06060606",
        398 => x"06060606",

                --  sprite 2
        399 => x"00010102",
        400 => x"02020202",
        401 => x"02020202",
        402 => x"02020200",
        403 => x"01000100",
        404 => x"00020200",
        405 => x"00000202",
        406 => x"01010101",
        407 => x"01010101",
        408 => x"01010101",
        409 => x"01010101",
        410 => x"01010101",
        411 => x"01000000",
        412 => x"00010101",
        413 => x"01010100",
        414 => x"00000002",
        415 => x"02020202",
        416 => x"00020202",
        417 => x"02020202",
        418 => x"02020202",
        419 => x"02020101",
        420 => x"02020201",
        421 => x"01010101",
        422 => x"01010101",
        423 => x"04010102",
        424 => x"02020202",
        425 => x"02020202",
        426 => x"02020204",
        427 => x"01040104",
        428 => x"04020204",
        429 => x"04040202",
        430 => x"01010101",
        431 => x"01010101",
        432 => x"01010101",
        433 => x"01010101",
        434 => x"01010101",
        435 => x"01040404",
        436 => x"04010101",
        437 => x"01010104",
        438 => x"04040402",
        439 => x"02020202",
        440 => x"04020202",
        441 => x"02020202",
        442 => x"02020202",
        443 => x"02020101",
        444 => x"02020201",
        445 => x"01010101",
        446 => x"01010101",
        447 => x"05060602",
        448 => x"02020202",
        449 => x"02020202",
        450 => x"02020205",
        451 => x"06050605",
        452 => x"05020205",
        453 => x"05050202",
        454 => x"06060606",
        455 => x"06060606",
        456 => x"06060606",
        457 => x"06060606",
        458 => x"06060606",
        459 => x"06050505",
        460 => x"05060606",
        461 => x"06060605",
        462 => x"05050502",
        463 => x"02020202",
        464 => x"05020202",
        465 => x"02020202",
        466 => x"02020202",
        467 => x"02020606",
        468 => x"02020206",
        469 => x"06060606",
        470 => x"06060606",

                --  sprite 3
        471 => x"00010100",
        472 => x"02020202",
        473 => x"02020202",
        474 => x"02020200",
        475 => x"00010000",
        476 => x"00020100",
        477 => x"00000000",
        478 => x"02010101",
        479 => x"01010101",
        480 => x"01010101",
        481 => x"01010101",
        482 => x"01010101",
        483 => x"01020000",
        484 => x"00010101",
        485 => x"01010100",
        486 => x"02000000",
        487 => x"00020202",
        488 => x"00020202",
        489 => x"02020202",
        490 => x"02020202",
        491 => x"02020202",
        492 => x"02020202",
        493 => x"01010101",
        494 => x"01010101",
        495 => x"04010104",
        496 => x"02020202",
        497 => x"02020202",
        498 => x"02020204",
        499 => x"04010404",
        500 => x"04020104",
        501 => x"04040404",
        502 => x"02010101",
        503 => x"01010101",
        504 => x"01010101",
        505 => x"01010101",
        506 => x"01010101",
        507 => x"01020404",
        508 => x"04010101",
        509 => x"01010104",
        510 => x"02040404",
        511 => x"04020202",
        512 => x"04020202",
        513 => x"02020202",
        514 => x"02020202",
        515 => x"02020202",
        516 => x"02020202",
        517 => x"01010101",
        518 => x"01010101",
        519 => x"05060605",
        520 => x"02020202",
        521 => x"02020202",
        522 => x"02020205",
        523 => x"05060505",
        524 => x"05020605",
        525 => x"05050505",
        526 => x"02060606",
        527 => x"06060606",
        528 => x"06060606",
        529 => x"06060606",
        530 => x"06060606",
        531 => x"06020505",
        532 => x"05060606",
        533 => x"06060605",
        534 => x"02050505",
        535 => x"05020202",
        536 => x"05020202",
        537 => x"02020202",
        538 => x"02020202",
        539 => x"02020202",
        540 => x"02020202",
        541 => x"06060606",
        542 => x"06060606",

                --  sprite 4
        543 => x"00010100",
        544 => x"01010102",
        545 => x"02020202",
        546 => x"02020200",
        547 => x"00010000",
        548 => x"00020100",
        549 => x"00000000",
        550 => x"02020101",
        551 => x"01010101",
        552 => x"01010101",
        553 => x"01010101",
        554 => x"01010101",
        555 => x"01030303",
        556 => x"00000001",
        557 => x"01010102",
        558 => x"02000000",
        559 => x"00000000",
        560 => x"00000202",
        561 => x"02020202",
        562 => x"02000000",
        563 => x"02020202",
        564 => x"02020202",
        565 => x"01010101",
        566 => x"01010101",
        567 => x"04010104",
        568 => x"01010102",
        569 => x"02020202",
        570 => x"02020204",
        571 => x"04010404",
        572 => x"04020104",
        573 => x"04040404",
        574 => x"02020101",
        575 => x"01010101",
        576 => x"01010101",
        577 => x"01010101",
        578 => x"01010101",
        579 => x"01030303",
        580 => x"04040401",
        581 => x"01010102",
        582 => x"02040404",
        583 => x"04040404",
        584 => x"04040202",
        585 => x"02020202",
        586 => x"02040404",
        587 => x"02020202",
        588 => x"02020202",
        589 => x"01010101",
        590 => x"01010101",
        591 => x"05060605",
        592 => x"06060602",
        593 => x"02020202",
        594 => x"02020205",
        595 => x"05060505",
        596 => x"05020605",
        597 => x"05050505",
        598 => x"02020606",
        599 => x"06060606",
        600 => x"06060606",
        601 => x"06060606",
        602 => x"06060606",
        603 => x"06030303",
        604 => x"05050506",
        605 => x"06060602",
        606 => x"02050505",
        607 => x"05050505",
        608 => x"05050202",
        609 => x"02020202",
        610 => x"02050505",
        611 => x"02020202",
        612 => x"02020202",
        613 => x"06060606",
        614 => x"06060606",

                --  sprite 5
        615 => x"00010100",
        616 => x"01010100",
        617 => x"02020202",
        618 => x"02020200",
        619 => x"00010000",
        620 => x"02010000",
        621 => x"00000000",
        622 => x"00020101",
        623 => x"01010101",
        624 => x"01010101",
        625 => x"01010101",
        626 => x"01010101",
        627 => x"03030303",
        628 => x"03000000",
        629 => x"01010102",
        630 => x"00000000",
        631 => x"00000000",
        632 => x"00000002",
        633 => x"02020200",
        634 => x"00000000",
        635 => x"02020202",
        636 => x"02000202",
        637 => x"01010101",
        638 => x"01010101",
        639 => x"04010104",
        640 => x"01010104",
        641 => x"02020202",
        642 => x"02020204",
        643 => x"04010404",
        644 => x"02010404",
        645 => x"04040404",
        646 => x"04020101",
        647 => x"01010101",
        648 => x"01010101",
        649 => x"01010101",
        650 => x"01010101",
        651 => x"03030303",
        652 => x"03040404",
        653 => x"01010102",
        654 => x"04040404",
        655 => x"04040404",
        656 => x"04040402",
        657 => x"02020204",
        658 => x"04040404",
        659 => x"02020202",
        660 => x"02040202",
        661 => x"01010101",
        662 => x"01010101",
        663 => x"05060605",
        664 => x"06060605",
        665 => x"02020202",
        666 => x"02020205",
        667 => x"05060505",
        668 => x"02060505",
        669 => x"05050505",
        670 => x"05020606",
        671 => x"06060606",
        672 => x"06060606",
        673 => x"06060606",
        674 => x"06060606",
        675 => x"03030303",
        676 => x"03050505",
        677 => x"06060602",
        678 => x"05050505",
        679 => x"05050505",
        680 => x"05050502",
        681 => x"02020205",
        682 => x"05050505",
        683 => x"02020202",
        684 => x"02050202",
        685 => x"06060606",
        686 => x"06060606",

                --  sprite 6
        687 => x"01020303",
        688 => x"03030303",
        689 => x"03030303",
        690 => x"03030102",
        691 => x"01010001",
        692 => x"00000000",
        693 => x"00020202",
        694 => x"02010101",
        695 => x"01010100",
        696 => x"00030202",
        697 => x"03000001",
        698 => x"01030101",
        699 => x"01010101",
        700 => x"01010101",
        701 => x"01010202",
        702 => x"00000200",
        703 => x"02020202",
        704 => x"02020202",
        705 => x"02020202",
        706 => x"02020202",
        707 => x"00020200",
        708 => x"02020002",
        709 => x"01010100",
        710 => x"00000201",
        711 => x"01020303",
        712 => x"03030303",
        713 => x"03030303",
        714 => x"03030102",
        715 => x"01010401",
        716 => x"04040404",
        717 => x"04020202",
        718 => x"02010101",
        719 => x"01010104",
        720 => x"04030202",
        721 => x"03040401",
        722 => x"01030101",
        723 => x"01010101",
        724 => x"01010101",
        725 => x"01010202",
        726 => x"04040204",
        727 => x"02020202",
        728 => x"02020202",
        729 => x"02020202",
        730 => x"02020202",
        731 => x"04020204",
        732 => x"02020402",
        733 => x"01010104",
        734 => x"04040201",
        735 => x"06020303",
        736 => x"03030303",
        737 => x"03030303",
        738 => x"03030602",
        739 => x"06060606",
        740 => x"05050505",
        741 => x"05050306",
        742 => x"06060606",
        743 => x"06060605",
        744 => x"05030202",
        745 => x"03050506",
        746 => x"06030606",
        747 => x"06060606",
        748 => x"06060606",
        749 => x"06060202",
        750 => x"05050205",
        751 => x"02020202",
        752 => x"02020202",
        753 => x"02020202",
        754 => x"02020202",
        755 => x"05020205",
        756 => x"02020502",
        757 => x"06060605",
        758 => x"05050206",

                --  sprite 7
        759 => x"01020303",
        760 => x"03030303",
        761 => x"03030303",
        762 => x"03030102",
        763 => x"01010000",
        764 => x"02000000",
        765 => x"00000202",
        766 => x"00020101",
        767 => x"01010100",
        768 => x"00030303",
        769 => x"03000001",
        770 => x"01030101",
        771 => x"01010101",
        772 => x"01010101",
        773 => x"01010002",
        774 => x"00000200",
        775 => x"02020202",
        776 => x"02020202",
        777 => x"02020202",
        778 => x"02020202",
        779 => x"00020200",
        780 => x"02020002",
        781 => x"01010002",
        782 => x"00020303",
        783 => x"01020303",
        784 => x"03030303",
        785 => x"03030303",
        786 => x"03030102",
        787 => x"01010404",
        788 => x"02040404",
        789 => x"04040202",
        790 => x"04020101",
        791 => x"01010104",
        792 => x"04030303",
        793 => x"03040401",
        794 => x"01030101",
        795 => x"01010101",
        796 => x"01010101",
        797 => x"01010402",
        798 => x"04040204",
        799 => x"02020202",
        800 => x"02020202",
        801 => x"02020202",
        802 => x"02020202",
        803 => x"04020204",
        804 => x"02020402",
        805 => x"01010402",
        806 => x"04020303",
        807 => x"06020303",
        808 => x"03030303",
        809 => x"03030303",
        810 => x"03030602",
        811 => x"06060605",
        812 => x"05050303",
        813 => x"02050503",
        814 => x"06060606",
        815 => x"06060605",
        816 => x"05030303",
        817 => x"03050506",
        818 => x"06030606",
        819 => x"06060606",
        820 => x"06060606",
        821 => x"06060502",
        822 => x"05050205",
        823 => x"02020202",
        824 => x"02020202",
        825 => x"02020202",
        826 => x"02020202",
        827 => x"05020205",
        828 => x"02020502",
        829 => x"06060502",
        830 => x"05020303",

                --  sprite 8
        831 => x"01020200",
        832 => x"00000000",
        833 => x"00000000",
        834 => x"00000102",
        835 => x"01000000",
        836 => x"00000000",
        837 => x"00000002",
        838 => x"02020101",
        839 => x"00000000",
        840 => x"00000200",
        841 => x"00000002",
        842 => x"01030101",
        843 => x"01010101",
        844 => x"01010101",
        845 => x"01010002",
        846 => x"00000200",
        847 => x"02020202",
        848 => x"02020202",
        849 => x"02020202",
        850 => x"02020202",
        851 => x"00020200",
        852 => x"00020202",
        853 => x"01000200",
        854 => x"02030301",
        855 => x"01020204",
        856 => x"04040404",
        857 => x"04040404",
        858 => x"04040102",
        859 => x"01040404",
        860 => x"04040404",
        861 => x"04040402",
        862 => x"02020101",
        863 => x"04040404",
        864 => x"04040204",
        865 => x"04040402",
        866 => x"01030101",
        867 => x"01010101",
        868 => x"01010101",
        869 => x"01010402",
        870 => x"04040204",
        871 => x"02020202",
        872 => x"02020202",
        873 => x"02020202",
        874 => x"02020202",
        875 => x"04020204",
        876 => x"04020202",
        877 => x"01040204",
        878 => x"02030301",
        879 => x"06020205",
        880 => x"05050505",
        881 => x"05050505",
        882 => x"05050602",
        883 => x"06060505",
        884 => x"05050303",
        885 => x"02050505",
        886 => x"03060606",
        887 => x"05050505",
        888 => x"05050205",
        889 => x"05050502",
        890 => x"06030606",
        891 => x"06060606",
        892 => x"06060606",
        893 => x"06060502",
        894 => x"05050205",
        895 => x"02020202",
        896 => x"02020202",
        897 => x"02020202",
        898 => x"02020202",
        899 => x"05020205",
        900 => x"05020202",
        901 => x"06050205",
        902 => x"02030306",

                --  sprite 9
        903 => x"01020303",
        904 => x"03030303",
        905 => x"03030303",
        906 => x"03030102",
        907 => x"01000000",
        908 => x"00000200",
        909 => x"00000200",
        910 => x"02020201",
        911 => x"00020000",
        912 => x"02000202",
        913 => x"02020200",
        914 => x"02030101",
        915 => x"01010101",
        916 => x"01010101",
        917 => x"01010002",
        918 => x"00000200",
        919 => x"02020202",
        920 => x"02020202",
        921 => x"02020202",
        922 => x"02020202",
        923 => x"00020200",
        924 => x"00000202",
        925 => x"00000202",
        926 => x"02010101",
        927 => x"01020303",
        928 => x"03030303",
        929 => x"03030303",
        930 => x"03030102",
        931 => x"01040404",
        932 => x"04040204",
        933 => x"04040204",
        934 => x"02020201",
        935 => x"04020404",
        936 => x"02040202",
        937 => x"02020204",
        938 => x"02030101",
        939 => x"01010101",
        940 => x"01010101",
        941 => x"01010402",
        942 => x"04040204",
        943 => x"02020202",
        944 => x"02020202",
        945 => x"02020202",
        946 => x"02020202",
        947 => x"04020204",
        948 => x"04040202",
        949 => x"04040202",
        950 => x"02010101",
        951 => x"06020303",
        952 => x"03030303",
        953 => x"03030303",
        954 => x"03030602",
        955 => x"06060505",
        956 => x"03030303",
        957 => x"03030205",
        958 => x"03060606",
        959 => x"05020505",
        960 => x"02050202",
        961 => x"02020205",
        962 => x"02030606",
        963 => x"06060606",
        964 => x"06060606",
        965 => x"06060502",
        966 => x"05050205",
        967 => x"02020202",
        968 => x"02020202",
        969 => x"02020202",
        970 => x"02020202",
        971 => x"05020205",
        972 => x"05050202",
        973 => x"05050202",
        974 => x"02060606",

                --  sprite 10
        975 => x"01020303",
        976 => x"03030303",
        977 => x"03030303",
        978 => x"03030102",
        979 => x"00000000",
        980 => x"00000000",
        981 => x"00000202",
        982 => x"02020101",
        983 => x"00000000",
        984 => x"00000200",
        985 => x"00000000",
        986 => x"00030201",
        987 => x"01010101",
        988 => x"01010101",
        989 => x"01010002",
        990 => x"00000200",
        991 => x"02020202",
        992 => x"02020202",
        993 => x"02020202",
        994 => x"02020202",
        995 => x"00020200",
        996 => x"02000200",
        997 => x"00020002",
        998 => x"01010101",
        999 => x"01020303",
        1000 => x"03030303",
        1001 => x"03030303",
        1002 => x"03030102",
        1003 => x"04040404",
        1004 => x"04040404",
        1005 => x"04040202",
        1006 => x"02020101",
        1007 => x"04040404",
        1008 => x"04040204",
        1009 => x"04040404",
        1010 => x"04030201",
        1011 => x"01010101",
        1012 => x"01010101",
        1013 => x"01010402",
        1014 => x"04040204",
        1015 => x"02020202",
        1016 => x"02020202",
        1017 => x"02020202",
        1018 => x"02020202",
        1019 => x"04020204",
        1020 => x"02040204",
        1021 => x"04020402",
        1022 => x"01010101",
        1023 => x"06020303",
        1024 => x"03030303",
        1025 => x"03030303",
        1026 => x"03030602",
        1027 => x"06060505",
        1028 => x"03030303",
        1029 => x"03030205",
        1030 => x"03060606",
        1031 => x"05050505",
        1032 => x"05050205",
        1033 => x"05050505",
        1034 => x"05030206",
        1035 => x"06060606",
        1036 => x"06060606",
        1037 => x"06060502",
        1038 => x"05050205",
        1039 => x"02020202",
        1040 => x"02020202",
        1041 => x"02020202",
        1042 => x"02020202",
        1043 => x"05020205",
        1044 => x"02050205",
        1045 => x"05020502",
        1046 => x"06060606",

                --  sprite 11
        1047 => x"01020303",
        1048 => x"03030303",
        1049 => x"03030303",
        1050 => x"03030102",
        1051 => x"00000200",
        1052 => x"00000000",
        1053 => x"00000002",
        1054 => x"02020201",
        1055 => x"00000000",
        1056 => x"00000200",
        1057 => x"00000002",
        1058 => x"00000201",
        1059 => x"01010101",
        1060 => x"01010101",
        1061 => x"01010002",
        1062 => x"00000200",
        1063 => x"02020202",
        1064 => x"02020202",
        1065 => x"02020202",
        1066 => x"02020202",
        1067 => x"00020200",
        1068 => x"02000200",
        1069 => x"02020002",
        1070 => x"01010101",
        1071 => x"01020303",
        1072 => x"03030303",
        1073 => x"03030303",
        1074 => x"03030102",
        1075 => x"04040204",
        1076 => x"04040404",
        1077 => x"04040402",
        1078 => x"02020201",
        1079 => x"04040404",
        1080 => x"04040204",
        1081 => x"04040402",
        1082 => x"04040201",
        1083 => x"01010101",
        1084 => x"01010101",
        1085 => x"01010402",
        1086 => x"04040204",
        1087 => x"02020202",
        1088 => x"02020202",
        1089 => x"02020202",
        1090 => x"02020202",
        1091 => x"04020204",
        1092 => x"02040204",
        1093 => x"02020402",
        1094 => x"01010101",
        1095 => x"06020303",
        1096 => x"03030303",
        1097 => x"03030303",
        1098 => x"03030602",
        1099 => x"06060505",
        1100 => x"02020303",
        1101 => x"02020205",
        1102 => x"03060606",
        1103 => x"05050505",
        1104 => x"05050205",
        1105 => x"05050502",
        1106 => x"05050206",
        1107 => x"06060606",
        1108 => x"06060606",
        1109 => x"06060502",
        1110 => x"05050205",
        1111 => x"02020202",
        1112 => x"02020202",
        1113 => x"02020202",
        1114 => x"02020202",
        1115 => x"05020205",
        1116 => x"02050205",
        1117 => x"02020502",
        1118 => x"06060606",

                --  sprite 12
        1119 => x"01010101",
        1120 => x"01010202",
        1121 => x"01000000",
        1122 => x"00000202",
        1123 => x"01000000",
        1124 => x"00000202",
        1125 => x"02000000",
        1126 => x"00000201",
        1127 => x"02000000",
        1128 => x"00000201",
        1129 => x"01010101",
        1130 => x"01010101",
        1131 => x"01010101",
        1132 => x"01010101",
        1133 => x"01010103",
        1134 => x"03000000",
        1135 => x"00030303",
        1136 => x"03030000",
        1137 => x"00000303",
        1138 => x"03030300",
        1139 => x"00000202",
        1140 => x"02010101",
        1141 => x"01010101",
        1142 => x"01010101",
        1143 => x"01010101",
        1144 => x"01010202",
        1145 => x"01040404",
        1146 => x"04040202",
        1147 => x"01040404",
        1148 => x"04040202",
        1149 => x"02040404",
        1150 => x"04040201",
        1151 => x"02040404",
        1152 => x"04040201",
        1153 => x"01010101",
        1154 => x"01010101",
        1155 => x"01010101",
        1156 => x"01010101",
        1157 => x"01010103",
        1158 => x"03040404",
        1159 => x"04030303",
        1160 => x"03030404",
        1161 => x"04040303",
        1162 => x"03030304",
        1163 => x"04040202",
        1164 => x"02010101",
        1165 => x"01010101",
        1166 => x"01010101",
        1167 => x"06060606",
        1168 => x"06060202",
        1169 => x"06050505",
        1170 => x"05050202",
        1171 => x"06050505",
        1172 => x"05050202",
        1173 => x"02050505",
        1174 => x"05050206",
        1175 => x"02050505",
        1176 => x"05050206",
        1177 => x"06060606",
        1178 => x"06060606",
        1179 => x"06060606",
        1180 => x"06060606",
        1181 => x"06060603",
        1182 => x"03050505",
        1183 => x"02060305",
        1184 => x"05030303",
        1185 => x"03030305",
        1186 => x"05020603",
        1187 => x"05050202",
        1188 => x"02060606",
        1189 => x"06060606",
        1190 => x"06060606",

                --  sprite 13
        1191 => x"01010101",
        1192 => x"01010002",
        1193 => x"01000000",
        1194 => x"00020202",
        1195 => x"01000000",
        1196 => x"00020202",
        1197 => x"01000000",
        1198 => x"00000002",
        1199 => x"01000000",
        1200 => x"00000002",
        1201 => x"01010101",
        1202 => x"01010101",
        1203 => x"01010101",
        1204 => x"01010101",
        1205 => x"01010300",
        1206 => x"00000000",
        1207 => x"03000000",
        1208 => x"00000200",
        1209 => x"00030000",
        1210 => x"00000002",
        1211 => x"00000000",
        1212 => x"02020101",
        1213 => x"01010101",
        1214 => x"01010101",
        1215 => x"01010101",
        1216 => x"01010402",
        1217 => x"01040404",
        1218 => x"04020202",
        1219 => x"01040404",
        1220 => x"04020202",
        1221 => x"01040404",
        1222 => x"04040402",
        1223 => x"01040404",
        1224 => x"04040402",
        1225 => x"01010101",
        1226 => x"01010101",
        1227 => x"01010101",
        1228 => x"01010101",
        1229 => x"01010304",
        1230 => x"04040404",
        1231 => x"03040404",
        1232 => x"04040204",
        1233 => x"04030404",
        1234 => x"04040402",
        1235 => x"04040404",
        1236 => x"02020101",
        1237 => x"01010101",
        1238 => x"01010101",
        1239 => x"06060606",
        1240 => x"06060502",
        1241 => x"06050505",
        1242 => x"05020202",
        1243 => x"06050505",
        1244 => x"05020202",
        1245 => x"06050505",
        1246 => x"05050502",
        1247 => x"06050505",
        1248 => x"05050502",
        1249 => x"06060606",
        1250 => x"06060606",
        1251 => x"06060606",
        1252 => x"06060606",
        1253 => x"06060305",
        1254 => x"05050505",
        1255 => x"05030505",
        1256 => x"03050202",
        1257 => x"02020502",
        1258 => x"05050205",
        1259 => x"05050505",
        1260 => x"02020606",
        1261 => x"06060606",
        1262 => x"06060606",

                --  sprite 14
        1263 => x"01010101",
        1264 => x"01000002",
        1265 => x"01000000",
        1266 => x"00000202",
        1267 => x"01000000",
        1268 => x"00000202",
        1269 => x"01000000",
        1270 => x"00000002",
        1271 => x"01000000",
        1272 => x"00000002",
        1273 => x"00010101",
        1274 => x"01010101",
        1275 => x"01010101",
        1276 => x"01010101",
        1277 => x"01010302",
        1278 => x"03000003",
        1279 => x"00000000",
        1280 => x"00000200",
        1281 => x"00030000",
        1282 => x"00000000",
        1283 => x"02000002",
        1284 => x"03020101",
        1285 => x"01010101",
        1286 => x"01010101",
        1287 => x"01010101",
        1288 => x"01040402",
        1289 => x"01040404",
        1290 => x"04040202",
        1291 => x"01040404",
        1292 => x"04040202",
        1293 => x"01040404",
        1294 => x"04040402",
        1295 => x"01040404",
        1296 => x"04040402",
        1297 => x"04010101",
        1298 => x"01010101",
        1299 => x"01010101",
        1300 => x"01010101",
        1301 => x"01010302",
        1302 => x"03040403",
        1303 => x"04040404",
        1304 => x"04040204",
        1305 => x"04030404",
        1306 => x"04040404",
        1307 => x"02040402",
        1308 => x"03020101",
        1309 => x"01010101",
        1310 => x"01010101",
        1311 => x"06060606",
        1312 => x"06050502",
        1313 => x"06050505",
        1314 => x"05050202",
        1315 => x"06050505",
        1316 => x"05050202",
        1317 => x"06050505",
        1318 => x"05050502",
        1319 => x"06050505",
        1320 => x"05050502",
        1321 => x"05060606",
        1322 => x"06060606",
        1323 => x"06060606",
        1324 => x"06060606",
        1325 => x"06060302",
        1326 => x"03050505",
        1327 => x"05050503",
        1328 => x"05050202",
        1329 => x"02020505",
        1330 => x"02050505",
        1331 => x"02050502",
        1332 => x"03020606",
        1333 => x"06060606",
        1334 => x"06060606",

                --  sprite 15
        1335 => x"01010101",
        1336 => x"01000002",
        1337 => x"02000000",
        1338 => x"00000201",
        1339 => x"02000000",
        1340 => x"00000201",
        1341 => x"01000000",
        1342 => x"00000202",
        1343 => x"01000000",
        1344 => x"00000202",
        1345 => x"00000202",
        1346 => x"02010101",
        1347 => x"01010101",
        1348 => x"01010101",
        1349 => x"01010302",
        1350 => x"03000003",
        1351 => x"02020202",
        1352 => x"02020200",
        1353 => x"00030202",
        1354 => x"02020202",
        1355 => x"02000002",
        1356 => x"03020101",
        1357 => x"01010101",
        1358 => x"01010101",
        1359 => x"01010101",
        1360 => x"01040402",
        1361 => x"02040404",
        1362 => x"04040201",
        1363 => x"02040404",
        1364 => x"04040201",
        1365 => x"01040404",
        1366 => x"04040202",
        1367 => x"01040404",
        1368 => x"04040202",
        1369 => x"04040202",
        1370 => x"02010101",
        1371 => x"01010101",
        1372 => x"01010101",
        1373 => x"01010302",
        1374 => x"03040403",
        1375 => x"02020202",
        1376 => x"02020204",
        1377 => x"04030202",
        1378 => x"02020202",
        1379 => x"02040402",
        1380 => x"03020101",
        1381 => x"01010101",
        1382 => x"01010101",
        1383 => x"06060606",
        1384 => x"06050502",
        1385 => x"02050505",
        1386 => x"05050206",
        1387 => x"02050505",
        1388 => x"05050206",
        1389 => x"06050505",
        1390 => x"05050202",
        1391 => x"06050505",
        1392 => x"05050202",
        1393 => x"05050202",
        1394 => x"02060606",
        1395 => x"06060606",
        1396 => x"06060606",
        1397 => x"06060302",
        1398 => x"03050505",
        1399 => x"05050503",
        1400 => x"05050505",
        1401 => x"05050505",
        1402 => x"02050505",
        1403 => x"02050502",
        1404 => x"03020606",
        1405 => x"06060606",
        1406 => x"06060606",

                --  sprite 16
        1407 => x"01010102",
        1408 => x"02000002",
        1409 => x"00000000",
        1410 => x"00000001",
        1411 => x"00000000",
        1412 => x"00000001",
        1413 => x"00000000",
        1414 => x"00000201",
        1415 => x"00000000",
        1416 => x"00000201",
        1417 => x"00020000",
        1418 => x"00020101",
        1419 => x"01010000",
        1420 => x"00000101",
        1421 => x"01010302",
        1422 => x"03000003",
        1423 => x"00000202",
        1424 => x"02000002",
        1425 => x"00030002",
        1426 => x"02020000",
        1427 => x"02000002",
        1428 => x"03020101",
        1429 => x"01010000",
        1430 => x"00000101",
        1431 => x"01010102",
        1432 => x"02040402",
        1433 => x"04040404",
        1434 => x"04040401",
        1435 => x"04040404",
        1436 => x"04040401",
        1437 => x"04040404",
        1438 => x"04040201",
        1439 => x"04040404",
        1440 => x"04040201",
        1441 => x"04020404",
        1442 => x"04020101",
        1443 => x"01010404",
        1444 => x"04040101",
        1445 => x"01010302",
        1446 => x"03040403",
        1447 => x"04040202",
        1448 => x"02040402",
        1449 => x"04030402",
        1450 => x"02020404",
        1451 => x"02040402",
        1452 => x"03020101",
        1453 => x"01010404",
        1454 => x"04040101",
        1455 => x"06060602",
        1456 => x"02050502",
        1457 => x"05050505",
        1458 => x"05050506",
        1459 => x"05050505",
        1460 => x"05050506",
        1461 => x"05050505",
        1462 => x"05050206",
        1463 => x"05050505",
        1464 => x"05050206",
        1465 => x"05020505",
        1466 => x"05020606",
        1467 => x"06060505",
        1468 => x"05050606",
        1469 => x"06060302",
        1470 => x"03050505",
        1471 => x"05050503",
        1472 => x"05050303",
        1473 => x"03030505",
        1474 => x"02050505",
        1475 => x"02050502",
        1476 => x"03020606",
        1477 => x"06060505",
        1478 => x"05050606",

                --  sprite 17
        1479 => x"01010000",
        1480 => x"02000002",
        1481 => x"00000000",
        1482 => x"00000001",
        1483 => x"00000000",
        1484 => x"00000001",
        1485 => x"00000000",
        1486 => x"00020201",
        1487 => x"00000000",
        1488 => x"00020201",
        1489 => x"00000000",
        1490 => x"00020101",
        1491 => x"01000000",
        1492 => x"00000001",
        1493 => x"01010302",
        1494 => x"03000003",
        1495 => x"00000000",
        1496 => x"00000002",
        1497 => x"00030000",
        1498 => x"00000000",
        1499 => x"02000002",
        1500 => x"03020101",
        1501 => x"01000000",
        1502 => x"00000001",
        1503 => x"01010404",
        1504 => x"02040402",
        1505 => x"04040404",
        1506 => x"04040401",
        1507 => x"04040404",
        1508 => x"04040401",
        1509 => x"04040404",
        1510 => x"04020201",
        1511 => x"04040404",
        1512 => x"04020201",
        1513 => x"04040404",
        1514 => x"04020101",
        1515 => x"01040404",
        1516 => x"04040401",
        1517 => x"01010302",
        1518 => x"03040403",
        1519 => x"04040404",
        1520 => x"04040402",
        1521 => x"04030404",
        1522 => x"04040404",
        1523 => x"02040402",
        1524 => x"03020101",
        1525 => x"01040404",
        1526 => x"04040401",
        1527 => x"06060505",
        1528 => x"02050502",
        1529 => x"05050505",
        1530 => x"05050506",
        1531 => x"05050505",
        1532 => x"05050506",
        1533 => x"05050505",
        1534 => x"05020206",
        1535 => x"05050505",
        1536 => x"05020206",
        1537 => x"05050505",
        1538 => x"05020606",
        1539 => x"06050505",
        1540 => x"05050506",
        1541 => x"06060302",
        1542 => x"03050505",
        1543 => x"05050505",
        1544 => x"02030205",
        1545 => x"05020302",
        1546 => x"05050505",
        1547 => x"02050502",
        1548 => x"03020606",
        1549 => x"06050505",
        1550 => x"05050506",

                --  sprite 18
        1551 => x"02000202",
        1552 => x"01000000",
        1553 => x"00000202",
        1554 => x"01000000",
        1555 => x"00000000",
        1556 => x"02010000",
        1557 => x"00000001",
        1558 => x"01020201",
        1559 => x"01000000",
        1560 => x"02000000",
        1561 => x"02020202",
        1562 => x"01010101",
        1563 => x"01010100",
        1564 => x"02010101",
        1565 => x"03020000",
        1566 => x"00000001",
        1567 => x"01010101",
        1568 => x"01010101",
        1569 => x"01010101",
        1570 => x"01010101",
        1571 => x"03000000",
        1572 => x"00020002",
        1573 => x"01010100",
        1574 => x"02010101",
        1575 => x"02040202",
        1576 => x"01040404",
        1577 => x"04040202",
        1578 => x"01040404",
        1579 => x"04040404",
        1580 => x"02010404",
        1581 => x"04040401",
        1582 => x"01020201",
        1583 => x"01040404",
        1584 => x"02040404",
        1585 => x"02020202",
        1586 => x"01010101",
        1587 => x"01010104",
        1588 => x"02010101",
        1589 => x"03020404",
        1590 => x"04040401",
        1591 => x"01010101",
        1592 => x"01010101",
        1593 => x"01010101",
        1594 => x"01010101",
        1595 => x"03040404",
        1596 => x"04020402",
        1597 => x"01010104",
        1598 => x"02010101",
        1599 => x"02050202",
        1600 => x"06050505",
        1601 => x"05050202",
        1602 => x"06050505",
        1603 => x"05050505",
        1604 => x"02060505",
        1605 => x"05050506",
        1606 => x"06020206",
        1607 => x"06050505",
        1608 => x"02050505",
        1609 => x"02020202",
        1610 => x"06060606",
        1611 => x"06060605",
        1612 => x"02060606",
        1613 => x"03020505",
        1614 => x"05050505",
        1615 => x"06060606",
        1616 => x"06060606",
        1617 => x"06060606",
        1618 => x"06060606",
        1619 => x"03050505",
        1620 => x"05020502",
        1621 => x"06060605",
        1622 => x"02060606",

                --  sprite 19
        1623 => x"01020202",
        1624 => x"01000000",
        1625 => x"00000202",
        1626 => x"02010000",
        1627 => x"00000000",
        1628 => x"02010000",
        1629 => x"00000100",
        1630 => x"00000201",
        1631 => x"01000000",
        1632 => x"02000000",
        1633 => x"02020101",
        1634 => x"01010101",
        1635 => x"01000000",
        1636 => x"00020201",
        1637 => x"03030202",
        1638 => x"02020201",
        1639 => x"01010101",
        1640 => x"00010101",
        1641 => x"01010101",
        1642 => x"01010101",
        1643 => x"02020202",
        1644 => x"02030002",
        1645 => x"01000000",
        1646 => x"00020201",
        1647 => x"01020202",
        1648 => x"01040404",
        1649 => x"04040202",
        1650 => x"02010404",
        1651 => x"04040404",
        1652 => x"02010404",
        1653 => x"04040104",
        1654 => x"04040201",
        1655 => x"01040404",
        1656 => x"02040404",
        1657 => x"02020101",
        1658 => x"01010101",
        1659 => x"01040404",
        1660 => x"04020201",
        1661 => x"03030202",
        1662 => x"02020201",
        1663 => x"01010101",
        1664 => x"04010101",
        1665 => x"01010101",
        1666 => x"01010101",
        1667 => x"02020202",
        1668 => x"02030402",
        1669 => x"01040404",
        1670 => x"04020201",
        1671 => x"06020202",
        1672 => x"06050505",
        1673 => x"05050202",
        1674 => x"02060505",
        1675 => x"05050505",
        1676 => x"02060505",
        1677 => x"05050605",
        1678 => x"05050206",
        1679 => x"06050505",
        1680 => x"02050505",
        1681 => x"02020606",
        1682 => x"06060606",
        1683 => x"06050505",
        1684 => x"05020206",
        1685 => x"03030202",
        1686 => x"02020205",
        1687 => x"06060606",
        1688 => x"05060606",
        1689 => x"06060606",
        1690 => x"06060606",
        1691 => x"02020202",
        1692 => x"02030502",
        1693 => x"06050505",
        1694 => x"05020206",

                --  sprite 20
        1695 => x"01010102",
        1696 => x"02000000",
        1697 => x"00000202",
        1698 => x"02010000",
        1699 => x"00000002",
        1700 => x"02010000",
        1701 => x"00000100",
        1702 => x"00000002",
        1703 => x"01000000",
        1704 => x"02000002",
        1705 => x"02010101",
        1706 => x"01010101",
        1707 => x"01030303",
        1708 => x"03030301",
        1709 => x"03020303",
        1710 => x"03030301",
        1711 => x"01010101",
        1712 => x"01010101",
        1713 => x"01010100",
        1714 => x"01010101",
        1715 => x"03030303",
        1716 => x"03000002",
        1717 => x"01030303",
        1718 => x"03030301",
        1719 => x"01010102",
        1720 => x"02040404",
        1721 => x"04040202",
        1722 => x"02010404",
        1723 => x"04040402",
        1724 => x"02010404",
        1725 => x"04040104",
        1726 => x"04040402",
        1727 => x"01040404",
        1728 => x"02040402",
        1729 => x"02010101",
        1730 => x"01010101",
        1731 => x"01030303",
        1732 => x"03030301",
        1733 => x"03020303",
        1734 => x"03030301",
        1735 => x"01010101",
        1736 => x"01010101",
        1737 => x"01010104",
        1738 => x"01010101",
        1739 => x"03030303",
        1740 => x"03040402",
        1741 => x"01030303",
        1742 => x"03030301",
        1743 => x"06060602",
        1744 => x"02050505",
        1745 => x"05050202",
        1746 => x"02060505",
        1747 => x"05050502",
        1748 => x"02060505",
        1749 => x"05050605",
        1750 => x"05050502",
        1751 => x"06050505",
        1752 => x"02050502",
        1753 => x"02060606",
        1754 => x"06060606",
        1755 => x"06030303",
        1756 => x"03030306",
        1757 => x"03020303",
        1758 => x"03030305",
        1759 => x"06060606",
        1760 => x"06060606",
        1761 => x"06060605",
        1762 => x"06060606",
        1763 => x"03030303",
        1764 => x"03050502",
        1765 => x"06030303",
        1766 => x"03030306",

                --  sprite 21
        1767 => x"01010101",
        1768 => x"02000200",
        1769 => x"00020202",
        1770 => x"02010000",
        1771 => x"00000002",
        1772 => x"02010000",
        1773 => x"00000100",
        1774 => x"00000002",
        1775 => x"01000000",
        1776 => x"02000002",
        1777 => x"02010101",
        1778 => x"01010101",
        1779 => x"03000000",
        1780 => x"00000002",
        1781 => x"03020000",
        1782 => x"00000001",
        1783 => x"01010101",
        1784 => x"01010100",
        1785 => x"01010101",
        1786 => x"01010101",
        1787 => x"03000000",
        1788 => x"00020002",
        1789 => x"03000000",
        1790 => x"00000002",
        1791 => x"01010101",
        1792 => x"02040204",
        1793 => x"04020202",
        1794 => x"02010404",
        1795 => x"04040402",
        1796 => x"02010404",
        1797 => x"04040104",
        1798 => x"04040402",
        1799 => x"01040404",
        1800 => x"02040402",
        1801 => x"02010101",
        1802 => x"01010101",
        1803 => x"03040404",
        1804 => x"04040402",
        1805 => x"03020404",
        1806 => x"04040401",
        1807 => x"01010101",
        1808 => x"01010104",
        1809 => x"01010101",
        1810 => x"01010101",
        1811 => x"03040404",
        1812 => x"04020402",
        1813 => x"03040404",
        1814 => x"04040402",
        1815 => x"06060606",
        1816 => x"02050205",
        1817 => x"05020202",
        1818 => x"02060505",
        1819 => x"05050502",
        1820 => x"02060505",
        1821 => x"05050605",
        1822 => x"05050502",
        1823 => x"06050505",
        1824 => x"02050502",
        1825 => x"02060606",
        1826 => x"06060606",
        1827 => x"03050505",
        1828 => x"05050502",
        1829 => x"03020505",
        1830 => x"05050505",
        1831 => x"06060606",
        1832 => x"06060605",
        1833 => x"06060606",
        1834 => x"06060606",
        1835 => x"03050505",
        1836 => x"05020502",
        1837 => x"03050505",
        1838 => x"05050502",

                --  sprite 22
        1839 => x"01010101",
        1840 => x"01020202",
        1841 => x"02020202",
        1842 => x"02010000",
        1843 => x"01000202",
        1844 => x"02010200",
        1845 => x"00020100",
        1846 => x"00000202",
        1847 => x"02010000",
        1848 => x"02000002",
        1849 => x"02010101",
        1850 => x"01010101",
        1851 => x"03000000",
        1852 => x"00000002",
        1853 => x"03020000",
        1854 => x"00000001",
        1855 => x"01010001",
        1856 => x"01010101",
        1857 => x"01010101",
        1858 => x"01010101",
        1859 => x"03000000",
        1860 => x"00020002",
        1861 => x"03000000",
        1862 => x"00000002",
        1863 => x"01010101",
        1864 => x"01020202",
        1865 => x"02020202",
        1866 => x"02010404",
        1867 => x"01040202",
        1868 => x"02010204",
        1869 => x"04020104",
        1870 => x"04040202",
        1871 => x"02010404",
        1872 => x"02040402",
        1873 => x"02010101",
        1874 => x"01010101",
        1875 => x"03040404",
        1876 => x"04040402",
        1877 => x"03020404",
        1878 => x"04040401",
        1879 => x"01010401",
        1880 => x"01010101",
        1881 => x"01010101",
        1882 => x"01010101",
        1883 => x"03040404",
        1884 => x"04020402",
        1885 => x"03040404",
        1886 => x"04040402",
        1887 => x"06060606",
        1888 => x"06020202",
        1889 => x"02020202",
        1890 => x"02060505",
        1891 => x"06050202",
        1892 => x"02060205",
        1893 => x"05020605",
        1894 => x"05050202",
        1895 => x"02060505",
        1896 => x"02050502",
        1897 => x"02060606",
        1898 => x"06060606",
        1899 => x"03050505",
        1900 => x"05050502",
        1901 => x"03020505",
        1902 => x"05050505",
        1903 => x"06060506",
        1904 => x"06060606",
        1905 => x"06060606",
        1906 => x"06060606",
        1907 => x"03050505",
        1908 => x"05020502",
        1909 => x"03050505",
        1910 => x"05050502",

                --  sprite 23
        1911 => x"01010101",
        1912 => x"01010101",
        1913 => x"02020202",
        1914 => x"02010000",
        1915 => x"01000201",
        1916 => x"01010202",
        1917 => x"00020100",
        1918 => x"00000201",
        1919 => x"02010000",
        1920 => x"02000002",
        1921 => x"02010101",
        1922 => x"01010101",
        1923 => x"03000000",
        1924 => x"00000002",
        1925 => x"03030202",
        1926 => x"02020201",
        1927 => x"01010101",
        1928 => x"01010101",
        1929 => x"01010101",
        1930 => x"01010001",
        1931 => x"02020202",
        1932 => x"02030002",
        1933 => x"03000000",
        1934 => x"00000002",
        1935 => x"01010101",
        1936 => x"01010101",
        1937 => x"02020202",
        1938 => x"02010404",
        1939 => x"01040201",
        1940 => x"01010202",
        1941 => x"04020104",
        1942 => x"04040201",
        1943 => x"02010404",
        1944 => x"02040402",
        1945 => x"02010101",
        1946 => x"01010101",
        1947 => x"03040404",
        1948 => x"04040402",
        1949 => x"03030202",
        1950 => x"02020201",
        1951 => x"01010101",
        1952 => x"01010101",
        1953 => x"01010101",
        1954 => x"01010401",
        1955 => x"02020202",
        1956 => x"02030402",
        1957 => x"03040404",
        1958 => x"04040402",
        1959 => x"06060606",
        1960 => x"06060606",
        1961 => x"02020202",
        1962 => x"02060505",
        1963 => x"06050206",
        1964 => x"06060202",
        1965 => x"05020605",
        1966 => x"05050206",
        1967 => x"02060505",
        1968 => x"02050502",
        1969 => x"02060606",
        1970 => x"06060606",
        1971 => x"03050505",
        1972 => x"05050502",
        1973 => x"03030202",
        1974 => x"02020205",
        1975 => x"06060606",
        1976 => x"06060606",
        1977 => x"06060606",
        1978 => x"06060506",
        1979 => x"02020202",
        1980 => x"02030502",
        1981 => x"03050505",
        1982 => x"05050502",

                --  sprite 24
        1983 => x"01010203",
        1984 => x"03000303",
        1985 => x"03030303",
        1986 => x"03030303",
        1987 => x"03030303",
        1988 => x"03030303",
        1989 => x"03030303",
        1990 => x"03030303",
        1991 => x"03030303",
        1992 => x"03030303",
        1993 => x"00030303",
        1994 => x"03030302",
        1995 => x"01010201",
        1996 => x"01000101",
        1997 => x"01010101",
        1998 => x"01010101",
        1999 => x"01010101",
        2000 => x"01010101",
        2001 => x"01010101",
        2002 => x"01010101",
        2003 => x"01010101",
        2004 => x"01010101",
        2005 => x"00010101",
        2006 => x"01010102",
        2007 => x"01010203",
        2008 => x"03040303",
        2009 => x"03030303",
        2010 => x"03030303",
        2011 => x"03030303",
        2012 => x"03030303",
        2013 => x"03030303",
        2014 => x"03030303",
        2015 => x"03030303",
        2016 => x"03030303",
        2017 => x"04030303",
        2018 => x"03030302",
        2019 => x"01010201",
        2020 => x"01040101",
        2021 => x"01010101",
        2022 => x"01010101",
        2023 => x"01010101",
        2024 => x"01010101",
        2025 => x"01010101",
        2026 => x"01010101",
        2027 => x"01010101",
        2028 => x"01010101",
        2029 => x"04010101",
        2030 => x"01010102",
        2031 => x"06060203",
        2032 => x"03050303",
        2033 => x"03030303",
        2034 => x"03030303",
        2035 => x"03030303",
        2036 => x"03030303",
        2037 => x"03030303",
        2038 => x"03030303",
        2039 => x"03030303",
        2040 => x"03030303",
        2041 => x"05030303",
        2042 => x"03030302",
        2043 => x"06060206",
        2044 => x"06050606",
        2045 => x"06060606",
        2046 => x"06060606",
        2047 => x"06060606",
        2048 => x"06060606",
        2049 => x"06060606",
        2050 => x"06060606",
        2051 => x"06060606",
        2052 => x"06060606",
        2053 => x"05060606",
        2054 => x"06060602",

                --  sprite 25
        2055 => x"01020203",
        2056 => x"03030303",
        2057 => x"03030303",
        2058 => x"03030303",
        2059 => x"03030303",
        2060 => x"03030303",
        2061 => x"03030303",
        2062 => x"03030303",
        2063 => x"03030303",
        2064 => x"03030303",
        2065 => x"03030303",
        2066 => x"00030302",
        2067 => x"01020201",
        2068 => x"01010101",
        2069 => x"01010101",
        2070 => x"01010101",
        2071 => x"01010101",
        2072 => x"01010101",
        2073 => x"01010101",
        2074 => x"01010101",
        2075 => x"01010101",
        2076 => x"01010101",
        2077 => x"01010101",
        2078 => x"00010102",
        2079 => x"01020203",
        2080 => x"03030303",
        2081 => x"03030303",
        2082 => x"03030303",
        2083 => x"03030303",
        2084 => x"03030303",
        2085 => x"03030303",
        2086 => x"03030303",
        2087 => x"03030303",
        2088 => x"03030303",
        2089 => x"03030303",
        2090 => x"04030302",
        2091 => x"01020201",
        2092 => x"01010101",
        2093 => x"01010101",
        2094 => x"01010101",
        2095 => x"01010101",
        2096 => x"01010101",
        2097 => x"01010101",
        2098 => x"01010101",
        2099 => x"01010101",
        2100 => x"01010101",
        2101 => x"01010101",
        2102 => x"04010102",
        2103 => x"06020203",
        2104 => x"03030303",
        2105 => x"03030303",
        2106 => x"03030303",
        2107 => x"03030303",
        2108 => x"03030303",
        2109 => x"03030303",
        2110 => x"03030303",
        2111 => x"03030303",
        2112 => x"03030303",
        2113 => x"03030303",
        2114 => x"05030302",
        2115 => x"06020206",
        2116 => x"06060606",
        2117 => x"06060606",
        2118 => x"06060606",
        2119 => x"06060606",
        2120 => x"06060606",
        2121 => x"06060606",
        2122 => x"06060606",
        2123 => x"06060606",
        2124 => x"06060606",
        2125 => x"06060606",
        2126 => x"05060602",

                --  sprite 26
        2127 => x"01020303",
        2128 => x"03030303",
        2129 => x"03030003",
        2130 => x"03030303",
        2131 => x"03030003",
        2132 => x"03030303",
        2133 => x"03030003",
        2134 => x"03030303",
        2135 => x"03030003",
        2136 => x"03030303",
        2137 => x"03030303",
        2138 => x"03030302",
        2139 => x"01020101",
        2140 => x"01010101",
        2141 => x"01010001",
        2142 => x"01010101",
        2143 => x"01010001",
        2144 => x"01010101",
        2145 => x"01010001",
        2146 => x"01010101",
        2147 => x"01010001",
        2148 => x"01010101",
        2149 => x"01010101",
        2150 => x"01010102",
        2151 => x"01020303",
        2152 => x"03030303",
        2153 => x"03030403",
        2154 => x"03030303",
        2155 => x"03030403",
        2156 => x"03030303",
        2157 => x"03030403",
        2158 => x"03030303",
        2159 => x"03030403",
        2160 => x"03030303",
        2161 => x"03030303",
        2162 => x"03030302",
        2163 => x"01020101",
        2164 => x"01010101",
        2165 => x"01010401",
        2166 => x"01010101",
        2167 => x"01010401",
        2168 => x"01010101",
        2169 => x"01010401",
        2170 => x"01010101",
        2171 => x"01010401",
        2172 => x"01010101",
        2173 => x"01010101",
        2174 => x"01010102",
        2175 => x"06020303",
        2176 => x"03030303",
        2177 => x"03030503",
        2178 => x"03030303",
        2179 => x"03030503",
        2180 => x"03030303",
        2181 => x"03030503",
        2182 => x"03030303",
        2183 => x"03030503",
        2184 => x"03030303",
        2185 => x"03030303",
        2186 => x"03030302",
        2187 => x"06020606",
        2188 => x"06060606",
        2189 => x"06060506",
        2190 => x"06060606",
        2191 => x"06060506",
        2192 => x"06060606",
        2193 => x"06060506",
        2194 => x"06060606",
        2195 => x"06060506",
        2196 => x"06060606",
        2197 => x"06060606",
        2198 => x"06060602",

                --  sprite 27
        2199 => x"01030300",
        2200 => x"03030303",
        2201 => x"03030303",
        2202 => x"03030303",
        2203 => x"03030303",
        2204 => x"03030303",
        2205 => x"03030303",
        2206 => x"03030303",
        2207 => x"03030303",
        2208 => x"03030303",
        2209 => x"03030303",
        2210 => x"03030301",
        2211 => x"01010100",
        2212 => x"01010101",
        2213 => x"01010101",
        2214 => x"01010101",
        2215 => x"01010101",
        2216 => x"01010101",
        2217 => x"01010101",
        2218 => x"01010101",
        2219 => x"01010101",
        2220 => x"01010101",
        2221 => x"01010101",
        2222 => x"01010101",
        2223 => x"01030304",
        2224 => x"03030303",
        2225 => x"03030303",
        2226 => x"03030303",
        2227 => x"03030303",
        2228 => x"03030303",
        2229 => x"03030303",
        2230 => x"03030303",
        2231 => x"03030303",
        2232 => x"03030303",
        2233 => x"03030303",
        2234 => x"03030301",
        2235 => x"01010104",
        2236 => x"01010101",
        2237 => x"01010101",
        2238 => x"01010101",
        2239 => x"01010101",
        2240 => x"01010101",
        2241 => x"01010101",
        2242 => x"01010101",
        2243 => x"01010101",
        2244 => x"01010101",
        2245 => x"01010101",
        2246 => x"01010101",
        2247 => x"06030305",
        2248 => x"03030303",
        2249 => x"03030303",
        2250 => x"03030303",
        2251 => x"03030303",
        2252 => x"03030303",
        2253 => x"03030303",
        2254 => x"03030303",
        2255 => x"03030303",
        2256 => x"03030303",
        2257 => x"03030303",
        2258 => x"03030306",
        2259 => x"06060605",
        2260 => x"06060606",
        2261 => x"06060606",
        2262 => x"06060606",
        2263 => x"06060606",
        2264 => x"06060606",
        2265 => x"06060606",
        2266 => x"06060606",
        2267 => x"06060606",
        2268 => x"06060606",
        2269 => x"06060606",
        2270 => x"06060606",

                --  sprite 28
        2271 => x"01030303",
        2272 => x"03030303",
        2273 => x"03030303",
        2274 => x"03030303",
        2275 => x"03030303",
        2276 => x"03030303",
        2277 => x"03030303",
        2278 => x"03030303",
        2279 => x"03030303",
        2280 => x"03030303",
        2281 => x"03030300",
        2282 => x"03030301",
        2283 => x"01010101",
        2284 => x"01010101",
        2285 => x"01010101",
        2286 => x"01010101",
        2287 => x"01010101",
        2288 => x"01010101",
        2289 => x"01010101",
        2290 => x"01010101",
        2291 => x"01010101",
        2292 => x"01010101",
        2293 => x"01010100",
        2294 => x"01010101",
        2295 => x"01030303",
        2296 => x"03030303",
        2297 => x"03030303",
        2298 => x"03030303",
        2299 => x"03030303",
        2300 => x"03030303",
        2301 => x"03030303",
        2302 => x"03030303",
        2303 => x"03030303",
        2304 => x"03030303",
        2305 => x"03030304",
        2306 => x"03030301",
        2307 => x"01010101",
        2308 => x"01010101",
        2309 => x"01010101",
        2310 => x"01010101",
        2311 => x"01010101",
        2312 => x"01010101",
        2313 => x"01010101",
        2314 => x"01010101",
        2315 => x"01010101",
        2316 => x"01010101",
        2317 => x"01010104",
        2318 => x"01010101",
        2319 => x"06030303",
        2320 => x"03030303",
        2321 => x"03030303",
        2322 => x"03030303",
        2323 => x"03030303",
        2324 => x"03030303",
        2325 => x"03030303",
        2326 => x"03030303",
        2327 => x"03030303",
        2328 => x"03030303",
        2329 => x"03030305",
        2330 => x"03030306",
        2331 => x"06060606",
        2332 => x"06060606",
        2333 => x"06060606",
        2334 => x"06060606",
        2335 => x"06060606",
        2336 => x"06060606",
        2337 => x"06060606",
        2338 => x"06060606",
        2339 => x"06060606",
        2340 => x"06060606",
        2341 => x"06060605",
        2342 => x"06060606",

                --  sprite 29
        2343 => x"01030303",
        2344 => x"03030003",
        2345 => x"03030303",
        2346 => x"03030303",
        2347 => x"03030303",
        2348 => x"03030303",
        2349 => x"03030303",
        2350 => x"03030303",
        2351 => x"03030303",
        2352 => x"03030303",
        2353 => x"03030303",
        2354 => x"03030101",
        2355 => x"01010101",
        2356 => x"01010001",
        2357 => x"01010101",
        2358 => x"01010101",
        2359 => x"01010101",
        2360 => x"01010101",
        2361 => x"01010101",
        2362 => x"01010101",
        2363 => x"01010101",
        2364 => x"01010101",
        2365 => x"01010101",
        2366 => x"01010101",
        2367 => x"01030303",
        2368 => x"03030403",
        2369 => x"03030303",
        2370 => x"03030303",
        2371 => x"03030303",
        2372 => x"03030303",
        2373 => x"03030303",
        2374 => x"03030303",
        2375 => x"03030303",
        2376 => x"03030303",
        2377 => x"03030303",
        2378 => x"03030101",
        2379 => x"01010101",
        2380 => x"01010401",
        2381 => x"01010101",
        2382 => x"01010101",
        2383 => x"01010101",
        2384 => x"01010101",
        2385 => x"01010101",
        2386 => x"01010101",
        2387 => x"01010101",
        2388 => x"01010101",
        2389 => x"01010101",
        2390 => x"01010101",
        2391 => x"06030303",
        2392 => x"03030503",
        2393 => x"03030303",
        2394 => x"03030303",
        2395 => x"03030303",
        2396 => x"03030303",
        2397 => x"03030303",
        2398 => x"03030303",
        2399 => x"03030303",
        2400 => x"03030303",
        2401 => x"03030303",
        2402 => x"03030606",
        2403 => x"06060606",
        2404 => x"06060506",
        2405 => x"06060606",
        2406 => x"06060606",
        2407 => x"06060606",
        2408 => x"06060606",
        2409 => x"06060606",
        2410 => x"06060606",
        2411 => x"06060606",
        2412 => x"06060606",
        2413 => x"06060606",
        2414 => x"06060606",

                --  sprite 30
        2415 => x"03030303",
        2416 => x"03030303",
        2417 => x"03030303",
        2418 => x"03030303",
        2419 => x"03030303",
        2420 => x"03030303",
        2421 => x"03030303",
        2422 => x"03030303",
        2423 => x"03030303",
        2424 => x"03030303",
        2425 => x"03030303",
        2426 => x"03030201",
        2427 => x"01010101",
        2428 => x"01010101",
        2429 => x"01010101",
        2430 => x"01010101",
        2431 => x"01010101",
        2432 => x"01010101",
        2433 => x"01010101",
        2434 => x"01010101",
        2435 => x"01010101",
        2436 => x"01010101",
        2437 => x"01010101",
        2438 => x"01010201",
        2439 => x"03030303",
        2440 => x"03030303",
        2441 => x"03030303",
        2442 => x"03030303",
        2443 => x"03030303",
        2444 => x"03030303",
        2445 => x"03030303",
        2446 => x"03030303",
        2447 => x"03030303",
        2448 => x"03030303",
        2449 => x"03030303",
        2450 => x"03030201",
        2451 => x"01010101",
        2452 => x"01010101",
        2453 => x"01010101",
        2454 => x"01010101",
        2455 => x"01010101",
        2456 => x"01010101",
        2457 => x"01010101",
        2458 => x"01010101",
        2459 => x"01010101",
        2460 => x"01010101",
        2461 => x"01010101",
        2462 => x"01010201",
        2463 => x"03030303",
        2464 => x"03030303",
        2465 => x"03030303",
        2466 => x"03030303",
        2467 => x"03030303",
        2468 => x"03030303",
        2469 => x"03030303",
        2470 => x"03030303",
        2471 => x"03030303",
        2472 => x"03030303",
        2473 => x"03030303",
        2474 => x"03030206",
        2475 => x"06060606",
        2476 => x"06060606",
        2477 => x"06060606",
        2478 => x"06060606",
        2479 => x"06060606",
        2480 => x"06060606",
        2481 => x"06060606",
        2482 => x"06060606",
        2483 => x"06060606",
        2484 => x"06060606",
        2485 => x"06060606",
        2486 => x"06060206",

                --  sprite 31
        2487 => x"03030303",
        2488 => x"03030303",
        2489 => x"03030303",
        2490 => x"03030303",
        2491 => x"03030303",
        2492 => x"03030303",
        2493 => x"03030303",
        2494 => x"03030303",
        2495 => x"03030303",
        2496 => x"03030303",
        2497 => x"03030303",
        2498 => x"03030201",
        2499 => x"01010101",
        2500 => x"01010101",
        2501 => x"01010101",
        2502 => x"01010101",
        2503 => x"01010101",
        2504 => x"01010101",
        2505 => x"01010101",
        2506 => x"01010101",
        2507 => x"01010101",
        2508 => x"01010101",
        2509 => x"01010101",
        2510 => x"01010201",
        2511 => x"03030303",
        2512 => x"03030303",
        2513 => x"03030303",
        2514 => x"03030303",
        2515 => x"03030303",
        2516 => x"03030303",
        2517 => x"03030303",
        2518 => x"03030303",
        2519 => x"03030303",
        2520 => x"03030303",
        2521 => x"03030303",
        2522 => x"03030201",
        2523 => x"01010101",
        2524 => x"01010101",
        2525 => x"01010101",
        2526 => x"01010101",
        2527 => x"01010101",
        2528 => x"01010101",
        2529 => x"01010101",
        2530 => x"01010101",
        2531 => x"01010101",
        2532 => x"01010101",
        2533 => x"01010101",
        2534 => x"01010201",
        2535 => x"03030303",
        2536 => x"03030303",
        2537 => x"03030303",
        2538 => x"03030303",
        2539 => x"03030303",
        2540 => x"03030303",
        2541 => x"03030303",
        2542 => x"03030303",
        2543 => x"03030303",
        2544 => x"03030303",
        2545 => x"03030303",
        2546 => x"03030206",
        2547 => x"06060606",
        2548 => x"06060606",
        2549 => x"06060606",
        2550 => x"06060606",
        2551 => x"06060606",
        2552 => x"06060606",
        2553 => x"06060606",
        2554 => x"06060606",
        2555 => x"06060606",
        2556 => x"06060606",
        2557 => x"06060606",
        2558 => x"06060206",

                --  sprite 32
        2559 => x"01030300",
        2560 => x"03030303",
        2561 => x"03030303",
        2562 => x"03030303",
        2563 => x"03030303",
        2564 => x"03030303",
        2565 => x"03030303",
        2566 => x"03030303",
        2567 => x"03030303",
        2568 => x"03030303",
        2569 => x"03030303",
        2570 => x"03030201",
        2571 => x"01010100",
        2572 => x"01010101",
        2573 => x"01010101",
        2574 => x"01010101",
        2575 => x"01010101",
        2576 => x"01010101",
        2577 => x"01010101",
        2578 => x"01010101",
        2579 => x"01010101",
        2580 => x"01010101",
        2581 => x"01010101",
        2582 => x"01010201",
        2583 => x"01030304",
        2584 => x"03030303",
        2585 => x"03030303",
        2586 => x"03030303",
        2587 => x"03030303",
        2588 => x"03030303",
        2589 => x"03030303",
        2590 => x"03030303",
        2591 => x"03030303",
        2592 => x"03030303",
        2593 => x"03030303",
        2594 => x"03030201",
        2595 => x"01010104",
        2596 => x"01010101",
        2597 => x"01010101",
        2598 => x"01010101",
        2599 => x"01010101",
        2600 => x"01010101",
        2601 => x"01010101",
        2602 => x"01010101",
        2603 => x"01010101",
        2604 => x"01010101",
        2605 => x"01010101",
        2606 => x"01010201",
        2607 => x"06030305",
        2608 => x"03030303",
        2609 => x"03030303",
        2610 => x"03030303",
        2611 => x"03030303",
        2612 => x"03030303",
        2613 => x"03030303",
        2614 => x"03030303",
        2615 => x"03030303",
        2616 => x"03030303",
        2617 => x"03030303",
        2618 => x"03030206",
        2619 => x"06060605",
        2620 => x"06060606",
        2621 => x"06060606",
        2622 => x"06060606",
        2623 => x"06060606",
        2624 => x"06060606",
        2625 => x"06060606",
        2626 => x"06060606",
        2627 => x"06060606",
        2628 => x"06060606",
        2629 => x"06060606",
        2630 => x"06060206",

                --  sprite 33
        2631 => x"01030303",
        2632 => x"03030303",
        2633 => x"03030300",
        2634 => x"03030303",
        2635 => x"03030300",
        2636 => x"03030303",
        2637 => x"03030300",
        2638 => x"03030303",
        2639 => x"03030300",
        2640 => x"03030303",
        2641 => x"03030300",
        2642 => x"03030201",
        2643 => x"01010101",
        2644 => x"01010101",
        2645 => x"01010100",
        2646 => x"01010101",
        2647 => x"01010100",
        2648 => x"01010101",
        2649 => x"01010100",
        2650 => x"01010101",
        2651 => x"01010100",
        2652 => x"01010101",
        2653 => x"01010100",
        2654 => x"01010201",
        2655 => x"01030303",
        2656 => x"03030303",
        2657 => x"03030304",
        2658 => x"03030303",
        2659 => x"03030304",
        2660 => x"03030303",
        2661 => x"03030304",
        2662 => x"03030303",
        2663 => x"03030304",
        2664 => x"03030303",
        2665 => x"03030304",
        2666 => x"03030201",
        2667 => x"01010101",
        2668 => x"01010101",
        2669 => x"01010104",
        2670 => x"01010101",
        2671 => x"01010104",
        2672 => x"01010101",
        2673 => x"01010104",
        2674 => x"01010101",
        2675 => x"01010104",
        2676 => x"01010101",
        2677 => x"01010104",
        2678 => x"01010201",
        2679 => x"06030303",
        2680 => x"03030303",
        2681 => x"03030305",
        2682 => x"03030303",
        2683 => x"03030305",
        2684 => x"03030303",
        2685 => x"03030305",
        2686 => x"03030303",
        2687 => x"03030305",
        2688 => x"03030303",
        2689 => x"03030305",
        2690 => x"03030206",
        2691 => x"06060606",
        2692 => x"06060606",
        2693 => x"06060605",
        2694 => x"06060606",
        2695 => x"06060605",
        2696 => x"06060606",
        2697 => x"06060605",
        2698 => x"06060606",
        2699 => x"06060605",
        2700 => x"06060606",
        2701 => x"06060605",
        2702 => x"06060206",

                --  sprite 34
        2703 => x"01030303",
        2704 => x"03030303",
        2705 => x"03030303",
        2706 => x"03030303",
        2707 => x"03030303",
        2708 => x"03030303",
        2709 => x"03030303",
        2710 => x"03030303",
        2711 => x"03030303",
        2712 => x"03030303",
        2713 => x"03030303",
        2714 => x"03030202",
        2715 => x"01010101",
        2716 => x"01010101",
        2717 => x"01010101",
        2718 => x"01010101",
        2719 => x"01010101",
        2720 => x"01010101",
        2721 => x"01010101",
        2722 => x"01010101",
        2723 => x"01010101",
        2724 => x"01010101",
        2725 => x"01010101",
        2726 => x"01010202",
        2727 => x"01030303",
        2728 => x"03030303",
        2729 => x"03030303",
        2730 => x"03030303",
        2731 => x"03030303",
        2732 => x"03030303",
        2733 => x"03030303",
        2734 => x"03030303",
        2735 => x"03030303",
        2736 => x"03030303",
        2737 => x"03030303",
        2738 => x"03030202",
        2739 => x"01010101",
        2740 => x"01010101",
        2741 => x"01010101",
        2742 => x"01010101",
        2743 => x"01010101",
        2744 => x"01010101",
        2745 => x"01010101",
        2746 => x"01010101",
        2747 => x"01010101",
        2748 => x"01010101",
        2749 => x"01010101",
        2750 => x"01010202",
        2751 => x"06030303",
        2752 => x"03030303",
        2753 => x"03030303",
        2754 => x"03030303",
        2755 => x"03030303",
        2756 => x"03030303",
        2757 => x"03030303",
        2758 => x"03030303",
        2759 => x"03030303",
        2760 => x"03030303",
        2761 => x"03030303",
        2762 => x"03030202",
        2763 => x"06060606",
        2764 => x"06060606",
        2765 => x"06060606",
        2766 => x"06060606",
        2767 => x"06060606",
        2768 => x"06060606",
        2769 => x"06060606",
        2770 => x"06060606",
        2771 => x"06060606",
        2772 => x"06060606",
        2773 => x"06060606",
        2774 => x"06060202",

                --  sprite 35
        2775 => x"01030303",
        2776 => x"03030303",
        2777 => x"03030303",
        2778 => x"03030303",
        2779 => x"03030303",
        2780 => x"03030303",
        2781 => x"03030303",
        2782 => x"03030303",
        2783 => x"03030303",
        2784 => x"03030303",
        2785 => x"03030303",
        2786 => x"03030302",
        2787 => x"01010101",
        2788 => x"01010101",
        2789 => x"01010101",
        2790 => x"01010101",
        2791 => x"01010101",
        2792 => x"01010101",
        2793 => x"01010101",
        2794 => x"01010101",
        2795 => x"01010101",
        2796 => x"01010101",
        2797 => x"01010101",
        2798 => x"01010102",
        2799 => x"01030303",
        2800 => x"03030303",
        2801 => x"03030303",
        2802 => x"03030303",
        2803 => x"03030303",
        2804 => x"03030303",
        2805 => x"03030303",
        2806 => x"03030303",
        2807 => x"03030303",
        2808 => x"03030303",
        2809 => x"03030303",
        2810 => x"03030302",
        2811 => x"01010101",
        2812 => x"01010101",
        2813 => x"01010101",
        2814 => x"01010101",
        2815 => x"01010101",
        2816 => x"01010101",
        2817 => x"01010101",
        2818 => x"01010101",
        2819 => x"01010101",
        2820 => x"01010101",
        2821 => x"01010101",
        2822 => x"01010102",
        2823 => x"06030303",
        2824 => x"03030303",
        2825 => x"03030303",
        2826 => x"03030303",
        2827 => x"03030303",
        2828 => x"03030303",
        2829 => x"03030303",
        2830 => x"03030303",
        2831 => x"03030303",
        2832 => x"03030303",
        2833 => x"03030303",
        2834 => x"03030302",
        2835 => x"06060606",
        2836 => x"06060606",
        2837 => x"06060606",
        2838 => x"06060606",
        2839 => x"06060606",
        2840 => x"06060606",
        2841 => x"06060606",
        2842 => x"06060606",
        2843 => x"06060606",
        2844 => x"06060606",
        2845 => x"06060606",
        2846 => x"06060602",

                --  sprite 36
        2847 => x"01010101",
        2848 => x"02030303",
        2849 => x"03030303",
        2850 => x"03030303",
        2851 => x"03030303",
        2852 => x"03030303",
        2853 => x"03030303",
        2854 => x"03030303",
        2855 => x"03030303",
        2856 => x"03030303",
        2857 => x"03030303",
        2858 => x"02010101",
        2859 => x"01010101",
        2860 => x"02010101",
        2861 => x"01010101",
        2862 => x"01010101",
        2863 => x"01010101",
        2864 => x"01010101",
        2865 => x"01010101",
        2866 => x"01010101",
        2867 => x"01010101",
        2868 => x"01010101",
        2869 => x"01010101",
        2870 => x"02010101",
        2871 => x"01010101",
        2872 => x"02030303",
        2873 => x"03030303",
        2874 => x"03030303",
        2875 => x"03030303",
        2876 => x"03030303",
        2877 => x"03030303",
        2878 => x"03030303",
        2879 => x"03030303",
        2880 => x"03030303",
        2881 => x"03030303",
        2882 => x"02010101",
        2883 => x"01010101",
        2884 => x"02010101",
        2885 => x"01010101",
        2886 => x"01010101",
        2887 => x"01010101",
        2888 => x"01010101",
        2889 => x"01010101",
        2890 => x"01010101",
        2891 => x"01010101",
        2892 => x"01010101",
        2893 => x"01010101",
        2894 => x"02010101",
        2895 => x"06060606",
        2896 => x"02030303",
        2897 => x"03030303",
        2898 => x"03030303",
        2899 => x"03030303",
        2900 => x"03030303",
        2901 => x"03030303",
        2902 => x"03030303",
        2903 => x"03030303",
        2904 => x"03030303",
        2905 => x"03030303",
        2906 => x"02060606",
        2907 => x"06060606",
        2908 => x"02060606",
        2909 => x"06060606",
        2910 => x"06060606",
        2911 => x"06060606",
        2912 => x"06060606",
        2913 => x"06060606",
        2914 => x"06060606",
        2915 => x"06060606",
        2916 => x"06060606",
        2917 => x"06060606",
        2918 => x"02060606",

                --  sprite 37
        2919 => x"01010102",
        2920 => x"02030303",
        2921 => x"03030303",
        2922 => x"03030303",
        2923 => x"03030303",
        2924 => x"03030303",
        2925 => x"03030303",
        2926 => x"03030303",
        2927 => x"03030303",
        2928 => x"03030303",
        2929 => x"00030303",
        2930 => x"02020101",
        2931 => x"01010102",
        2932 => x"02010101",
        2933 => x"01010101",
        2934 => x"01010101",
        2935 => x"01010101",
        2936 => x"01010101",
        2937 => x"01010101",
        2938 => x"01010101",
        2939 => x"01010101",
        2940 => x"01010101",
        2941 => x"00010101",
        2942 => x"02020101",
        2943 => x"01010102",
        2944 => x"02030303",
        2945 => x"03030303",
        2946 => x"03030303",
        2947 => x"03030303",
        2948 => x"03030303",
        2949 => x"03030303",
        2950 => x"03030303",
        2951 => x"03030303",
        2952 => x"03030303",
        2953 => x"04030303",
        2954 => x"02020101",
        2955 => x"01010102",
        2956 => x"02010101",
        2957 => x"01010101",
        2958 => x"01010101",
        2959 => x"01010101",
        2960 => x"01010101",
        2961 => x"01010101",
        2962 => x"01010101",
        2963 => x"01010101",
        2964 => x"01010101",
        2965 => x"04010101",
        2966 => x"02020101",
        2967 => x"06060602",
        2968 => x"02030303",
        2969 => x"03030303",
        2970 => x"03030303",
        2971 => x"03030303",
        2972 => x"03030303",
        2973 => x"03030303",
        2974 => x"03030303",
        2975 => x"03030303",
        2976 => x"03030303",
        2977 => x"05030303",
        2978 => x"02020606",
        2979 => x"06060602",
        2980 => x"02060606",
        2981 => x"06060606",
        2982 => x"06060606",
        2983 => x"06060606",
        2984 => x"06060606",
        2985 => x"06060606",
        2986 => x"06060606",
        2987 => x"06060606",
        2988 => x"06060606",
        2989 => x"05060606",
        2990 => x"02020606",

                --  sprite 38
        2991 => x"01010101",
        2992 => x"01010303",
        2993 => x"00030300",
        2994 => x"03010303",
        2995 => x"00030300",
        2996 => x"03010303",
        2997 => x"00030300",
        2998 => x"03010303",
        2999 => x"00030300",
        3000 => x"03010303",
        3001 => x"03030301",
        3002 => x"01010101",
        3003 => x"01010101",
        3004 => x"01010101",
        3005 => x"00010100",
        3006 => x"01010101",
        3007 => x"00010100",
        3008 => x"01010101",
        3009 => x"00010100",
        3010 => x"01010101",
        3011 => x"00010100",
        3012 => x"01010101",
        3013 => x"01010101",
        3014 => x"01010101",
        3015 => x"01010101",
        3016 => x"01010303",
        3017 => x"04030304",
        3018 => x"03010303",
        3019 => x"04030304",
        3020 => x"03010303",
        3021 => x"04030304",
        3022 => x"03010303",
        3023 => x"04030304",
        3024 => x"03010303",
        3025 => x"03030301",
        3026 => x"01010101",
        3027 => x"01010101",
        3028 => x"01010101",
        3029 => x"04010104",
        3030 => x"01010101",
        3031 => x"04010104",
        3032 => x"01010101",
        3033 => x"04010104",
        3034 => x"01010101",
        3035 => x"04010104",
        3036 => x"01010101",
        3037 => x"01010101",
        3038 => x"01010101",
        3039 => x"06060606",
        3040 => x"06060303",
        3041 => x"05030305",
        3042 => x"03060303",
        3043 => x"05030305",
        3044 => x"03060303",
        3045 => x"05030305",
        3046 => x"03060303",
        3047 => x"05030305",
        3048 => x"03060303",
        3049 => x"03030306",
        3050 => x"06060606",
        3051 => x"06060606",
        3052 => x"06060606",
        3053 => x"05060605",
        3054 => x"06060606",
        3055 => x"05060605",
        3056 => x"06060606",
        3057 => x"05060605",
        3058 => x"06060606",
        3059 => x"05060605",
        3060 => x"06060606",
        3061 => x"06060606",
        3062 => x"06060606",

                --  sprite 39
        3063 => x"01010101",
        3064 => x"01010101",
        3065 => x"03030103",
        3066 => x"01010101",
        3067 => x"03030103",
        3068 => x"01010101",
        3069 => x"03030103",
        3070 => x"01010101",
        3071 => x"03030103",
        3072 => x"01010101",
        3073 => x"01010101",
        3074 => x"01010101",
        3075 => x"01010101",
        3076 => x"01010101",
        3077 => x"01010101",
        3078 => x"01010101",
        3079 => x"01010101",
        3080 => x"01010101",
        3081 => x"01010101",
        3082 => x"01010101",
        3083 => x"01010101",
        3084 => x"01010101",
        3085 => x"01010101",
        3086 => x"01010101",
        3087 => x"01010101",
        3088 => x"01010101",
        3089 => x"03030103",
        3090 => x"01010101",
        3091 => x"03030103",
        3092 => x"01010101",
        3093 => x"03030103",
        3094 => x"01010101",
        3095 => x"03030103",
        3096 => x"01010101",
        3097 => x"01010101",
        3098 => x"01010101",
        3099 => x"01010101",
        3100 => x"01010101",
        3101 => x"01010101",
        3102 => x"01010101",
        3103 => x"01010101",
        3104 => x"01010101",
        3105 => x"01010101",
        3106 => x"01010101",
        3107 => x"01010101",
        3108 => x"01010101",
        3109 => x"01010101",
        3110 => x"01010101",
        3111 => x"06060606",
        3112 => x"06060606",
        3113 => x"03030603",
        3114 => x"06060606",
        3115 => x"03030603",
        3116 => x"06060606",
        3117 => x"03030603",
        3118 => x"06060606",
        3119 => x"03030603",
        3120 => x"06060606",
        3121 => x"06060606",
        3122 => x"06060606",
        3123 => x"06060606",
        3124 => x"06060606",
        3125 => x"06060606",
        3126 => x"06060606",
        3127 => x"06060606",
        3128 => x"06060606",
        3129 => x"06060606",
        3130 => x"06060606",
        3131 => x"06060606",
        3132 => x"06060606",
        3133 => x"06060606",
        3134 => x"06060606",

                --  sprite 40
        3135 => x"03030300",
        3136 => x"03030303",
        3137 => x"01010101",
        3138 => x"01010101",
        3139 => x"01010101",
        3140 => x"01010101",
        3141 => x"03030303",
        3142 => x"03000303",
        3143 => x"01010101",
        3144 => x"01010101",
        3145 => x"01010101",
        3146 => x"01010101",
        3147 => x"01010101",
        3148 => x"01010101",
        3149 => x"01010101",
        3150 => x"01010101",
        3151 => x"03010303",
        3152 => x"03030303",
        3153 => x"00030302",
        3154 => x"03030303",
        3155 => x"00000000",
        3156 => x"00000003",
        3157 => x"00000000",
        3158 => x"00000003",
        3159 => x"03030304",
        3160 => x"03030303",
        3161 => x"01010101",
        3162 => x"01010101",
        3163 => x"01010101",
        3164 => x"01010101",
        3165 => x"03030303",
        3166 => x"03040303",
        3167 => x"01010101",
        3168 => x"01010101",
        3169 => x"01010101",
        3170 => x"01010101",
        3171 => x"01010101",
        3172 => x"01010101",
        3173 => x"01010101",
        3174 => x"01010101",
        3175 => x"03010303",
        3176 => x"03030303",
        3177 => x"04030302",
        3178 => x"03030303",
        3179 => x"04040404",
        3180 => x"04040403",
        3181 => x"04040404",
        3182 => x"04040403",
        3183 => x"03030305",
        3184 => x"03030303",
        3185 => x"06060606",
        3186 => x"06060606",
        3187 => x"06060606",
        3188 => x"06060606",
        3189 => x"03030303",
        3190 => x"03050303",
        3191 => x"06060606",
        3192 => x"06060606",
        3193 => x"06060606",
        3194 => x"06060606",
        3195 => x"06060606",
        3196 => x"06060606",
        3197 => x"06060606",
        3198 => x"06060606",
        3199 => x"03060303",
        3200 => x"03030303",
        3201 => x"05030302",
        3202 => x"03030303",
        3203 => x"05050505",
        3204 => x"05050503",
        3205 => x"05050505",
        3206 => x"05050503",

                --  sprite 41
        3207 => x"03030303",
        3208 => x"03030101",
        3209 => x"01010101",
        3210 => x"01010101",
        3211 => x"01010101",
        3212 => x"01010101",
        3213 => x"01030101",
        3214 => x"03030303",
        3215 => x"01010101",
        3216 => x"01010101",
        3217 => x"01010101",
        3218 => x"01010101",
        3219 => x"01010101",
        3220 => x"01010101",
        3221 => x"01010101",
        3222 => x"01010101",
        3223 => x"03010303",
        3224 => x"03020303",
        3225 => x"00030302",
        3226 => x"03000303",
        3227 => x"00020000",
        3228 => x"00020002",
        3229 => x"00020000",
        3230 => x"00020002",
        3231 => x"03030303",
        3232 => x"03030101",
        3233 => x"01010101",
        3234 => x"01010101",
        3235 => x"01010101",
        3236 => x"01010101",
        3237 => x"01030101",
        3238 => x"03030303",
        3239 => x"01010101",
        3240 => x"01010101",
        3241 => x"01010101",
        3242 => x"01010101",
        3243 => x"01010101",
        3244 => x"01010101",
        3245 => x"01010101",
        3246 => x"01010101",
        3247 => x"03010303",
        3248 => x"03020303",
        3249 => x"04030302",
        3250 => x"03040303",
        3251 => x"04020404",
        3252 => x"04020402",
        3253 => x"04020404",
        3254 => x"04020402",
        3255 => x"03030303",
        3256 => x"03030606",
        3257 => x"06060606",
        3258 => x"06060606",
        3259 => x"06060606",
        3260 => x"06060606",
        3261 => x"06030606",
        3262 => x"03030303",
        3263 => x"06060606",
        3264 => x"06060606",
        3265 => x"06060606",
        3266 => x"06060606",
        3267 => x"06060606",
        3268 => x"06060606",
        3269 => x"06060606",
        3270 => x"06060606",
        3271 => x"03060303",
        3272 => x"03020303",
        3273 => x"05030302",
        3274 => x"03050303",
        3275 => x"05020505",
        3276 => x"05020502",
        3277 => x"05020505",
        3278 => x"05020502",

                --  sprite 42
        3279 => x"01010101",
        3280 => x"01010101",
        3281 => x"01010101",
        3282 => x"01010101",
        3283 => x"01010101",
        3284 => x"01010101",
        3285 => x"01010101",
        3286 => x"01010101",
        3287 => x"03000302",
        3288 => x"02020201",
        3289 => x"01010101",
        3290 => x"01010101",
        3291 => x"01010101",
        3292 => x"01010101",
        3293 => x"01010102",
        3294 => x"02030303",
        3295 => x"03030303",
        3296 => x"03030303",
        3297 => x"03030303",
        3298 => x"03030303",
        3299 => x"00000000",
        3300 => x"00000002",
        3301 => x"00000000",
        3302 => x"00000002",
        3303 => x"01010101",
        3304 => x"01010101",
        3305 => x"01010101",
        3306 => x"01010101",
        3307 => x"01010101",
        3308 => x"01010101",
        3309 => x"01010101",
        3310 => x"01010101",
        3311 => x"03040302",
        3312 => x"02020201",
        3313 => x"01010101",
        3314 => x"01010101",
        3315 => x"01010101",
        3316 => x"01010101",
        3317 => x"01010102",
        3318 => x"02030303",
        3319 => x"03030303",
        3320 => x"03030303",
        3321 => x"03030303",
        3322 => x"03030303",
        3323 => x"04040404",
        3324 => x"04040402",
        3325 => x"04040404",
        3326 => x"04040402",
        3327 => x"06060606",
        3328 => x"06060606",
        3329 => x"06060606",
        3330 => x"06060606",
        3331 => x"06060606",
        3332 => x"06060606",
        3333 => x"06060606",
        3334 => x"06060606",
        3335 => x"03050302",
        3336 => x"02020206",
        3337 => x"06060606",
        3338 => x"06060606",
        3339 => x"06060606",
        3340 => x"06060606",
        3341 => x"06060602",
        3342 => x"02030303",
        3343 => x"03030303",
        3344 => x"03030303",
        3345 => x"03030303",
        3346 => x"03030303",
        3347 => x"05050505",
        3348 => x"05050502",
        3349 => x"05050505",
        3350 => x"05050502",

                --  sprite 43
        3351 => x"01010101",
        3352 => x"01010101",
        3353 => x"01010101",
        3354 => x"01010101",
        3355 => x"01010101",
        3356 => x"01010101",
        3357 => x"01010101",
        3358 => x"01010101",
        3359 => x"03030303",
        3360 => x"03030202",
        3361 => x"01010101",
        3362 => x"01010101",
        3363 => x"01010101",
        3364 => x"01010101",
        3365 => x"02020203",
        3366 => x"03030300",
        3367 => x"03030303",
        3368 => x"03030303",
        3369 => x"03030303",
        3370 => x"03030303",
        3371 => x"03020202",
        3372 => x"02020202",
        3373 => x"03020202",
        3374 => x"02020202",
        3375 => x"01010101",
        3376 => x"01010101",
        3377 => x"01010101",
        3378 => x"01010101",
        3379 => x"01010101",
        3380 => x"01010101",
        3381 => x"01010101",
        3382 => x"01010101",
        3383 => x"03030303",
        3384 => x"03030202",
        3385 => x"01010101",
        3386 => x"01010101",
        3387 => x"01010101",
        3388 => x"01010101",
        3389 => x"02020203",
        3390 => x"03030304",
        3391 => x"03030303",
        3392 => x"03030303",
        3393 => x"03030303",
        3394 => x"03030303",
        3395 => x"03020202",
        3396 => x"02020202",
        3397 => x"03020202",
        3398 => x"02020202",
        3399 => x"06060606",
        3400 => x"06060606",
        3401 => x"06060606",
        3402 => x"06060606",
        3403 => x"06060606",
        3404 => x"06060606",
        3405 => x"06060606",
        3406 => x"06060606",
        3407 => x"03030303",
        3408 => x"03030202",
        3409 => x"06060606",
        3410 => x"06060606",
        3411 => x"06060606",
        3412 => x"06060606",
        3413 => x"02020203",
        3414 => x"03030307",
        3415 => x"03030303",
        3416 => x"03030303",
        3417 => x"03030303",
        3418 => x"03030303",
        3419 => x"03020202",
        3420 => x"02020202",
        3421 => x"03020202",
        3422 => x"02020202",

                --  sprite 44
        3423 => x"01010101",
        3424 => x"01010101",
        3425 => x"01010101",
        3426 => x"01010101",
        3427 => x"03010303",
        3428 => x"03030303",
        3429 => x"00030302",
        3430 => x"03030303",
        3431 => x"06060606",
        3432 => x"06060606",
        3433 => x"06060606",
        3434 => x"06060606",
        3435 => x"01010101",
        3436 => x"01010101",
        3437 => x"01010101",
        3438 => x"01010101",
        3439 => x"06060606",
        3440 => x"06060606",
        3441 => x"06060606",
        3442 => x"06060606",
        3443 => x"01010101",
        3444 => x"01010101",
        3445 => x"01010101",
        3446 => x"01010101",
        3447 => x"06060606",
        3448 => x"06030303",
        3449 => x"03030306",
        3450 => x"06060606",
        3451 => x"05050505",
        3452 => x"05050505",
        3453 => x"03050505",
        3454 => x"05050506",
        3455 => x"03050305",
        3456 => x"02050502",
        3457 => x"05050505",
        3458 => x"05050505",
        3459 => x"01010101",
        3460 => x"01010101",
        3461 => x"01010101",
        3462 => x"01010101",
        3463 => x"02020202",
        3464 => x"02020202",
        3465 => x"02020202",
        3466 => x"02020202",
        3467 => x"02020202",
        3468 => x"02020202",
        3469 => x"02020202",
        3470 => x"02020202",
        3471 => x"02020202",
        3472 => x"02020202",
        3473 => x"02020202",
        3474 => x"02020202",
        3475 => x"02020202",
        3476 => x"02020202",
        3477 => x"02020202",
        3478 => x"02020202",
        3479 => x"02020202",
        3480 => x"02020202",
        3481 => x"02020202",
        3482 => x"02020202",
        3483 => x"02020202",
        3484 => x"02020202",
        3485 => x"02020202",
        3486 => x"02020202",
        3487 => x"02020202",
        3488 => x"02020202",
        3489 => x"02020202",
        3490 => x"02020202",
        3491 => x"02020202",
        3492 => x"02020202",
        3493 => x"02020202",
        3494 => x"02020202",

                --  sprite 45
        3495 => x"01010101",
        3496 => x"01030303",
        3497 => x"03030301",
        3498 => x"01010103",
        3499 => x"03010303",
        3500 => x"03020303",
        3501 => x"00030302",
        3502 => x"03000303",
        3503 => x"06060606",
        3504 => x"05060502",
        3505 => x"02020606",
        3506 => x"06060606",
        3507 => x"01010101",
        3508 => x"00010002",
        3509 => x"02020101",
        3510 => x"01010101",
        3511 => x"06060606",
        3512 => x"06060606",
        3513 => x"06060606",
        3514 => x"06060303",
        3515 => x"01010101",
        3516 => x"04010402",
        3517 => x"02020101",
        3518 => x"01010101",
        3519 => x"03030303",
        3520 => x"03030505",
        3521 => x"05050503",
        3522 => x"03030303",
        3523 => x"02020202",
        3524 => x"02020202",
        3525 => x"03050505",
        3526 => x"05050506",
        3527 => x"03050305",
        3528 => x"02050502",
        3529 => x"02020202",
        3530 => x"02020202",
        3531 => x"01010101",
        3532 => x"01030303",
        3533 => x"03030301",
        3534 => x"01010103",
        3535 => x"02020202",
        3536 => x"02020202",
        3537 => x"02020202",
        3538 => x"02020202",
        3539 => x"02020202",
        3540 => x"02020202",
        3541 => x"02020202",
        3542 => x"02020202",
        3543 => x"02020202",
        3544 => x"02020202",
        3545 => x"02020202",
        3546 => x"02020202",
        3547 => x"02020202",
        3548 => x"02020202",
        3549 => x"02020202",
        3550 => x"02020202",
        3551 => x"02020202",
        3552 => x"02020202",
        3553 => x"02020202",
        3554 => x"02020202",
        3555 => x"02020202",
        3556 => x"02020202",
        3557 => x"02020202",
        3558 => x"02020202",
        3559 => x"02020202",
        3560 => x"02020202",
        3561 => x"02020202",
        3562 => x"02020202",
        3563 => x"02020202",
        3564 => x"02020202",
        3565 => x"02020202",
        3566 => x"02020202",

                --  sprite 46
        3567 => x"02010103",
        3568 => x"03000000",
        3569 => x"00000002",
        3570 => x"02010103",
        3571 => x"01010303",
        3572 => x"01020303",
        3573 => x"00000303",
        3574 => x"03000301",
        3575 => x"06060506",
        3576 => x"05050505",
        3577 => x"05020202",
        3578 => x"02060606",
        3579 => x"01010001",
        3580 => x"00000000",
        3581 => x"00020202",
        3582 => x"02010101",
        3583 => x"06060606",
        3584 => x"06060606",
        3585 => x"06060606",
        3586 => x"06030505",
        3587 => x"01010401",
        3588 => x"04040404",
        3589 => x"04020202",
        3590 => x"02010101",
        3591 => x"05050505",
        3592 => x"05020505",
        3593 => x"05050502",
        3594 => x"05050505",
        3595 => x"06050505",
        3596 => x"05050206",
        3597 => x"03020505",
        3598 => x"05050506",
        3599 => x"03050305",
        3600 => x"02020502",
        3601 => x"06050505",
        3602 => x"05050206",
        3603 => x"02010103",
        3604 => x"03040404",
        3605 => x"04040402",
        3606 => x"02010103",
        3607 => x"02020202",
        3608 => x"02020202",
        3609 => x"02020202",
        3610 => x"02020202",
        3611 => x"02020202",
        3612 => x"02020202",
        3613 => x"02020202",
        3614 => x"02020202",
        3615 => x"02020202",
        3616 => x"02020202",
        3617 => x"02020202",
        3618 => x"02020202",
        3619 => x"02020202",
        3620 => x"02020202",
        3621 => x"02020202",
        3622 => x"02020202",
        3623 => x"02020202",
        3624 => x"02020202",
        3625 => x"02020202",
        3626 => x"02020202",
        3627 => x"02020202",
        3628 => x"02020202",
        3629 => x"02020202",
        3630 => x"02020202",
        3631 => x"02020202",
        3632 => x"02020202",
        3633 => x"02020202",
        3634 => x"02020202",
        3635 => x"02020202",
        3636 => x"02020202",
        3637 => x"02020202",
        3638 => x"02020202",

                --  sprite 47
        3639 => x"02010300",
        3640 => x"00000000",
        3641 => x"00000000",
        3642 => x"00020103",
        3643 => x"00000303",
        3644 => x"01030103",
        3645 => x"00010300",
        3646 => x"03010101",
        3647 => x"06060505",
        3648 => x"02050505",
        3649 => x"05050202",
        3650 => x"05020606",
        3651 => x"01010000",
        3652 => x"02000000",
        3653 => x"00000202",
        3654 => x"00020101",
        3655 => x"06060606",
        3656 => x"06060606",
        3657 => x"06060606",
        3658 => x"06030505",
        3659 => x"01010404",
        3660 => x"02040404",
        3661 => x"04040202",
        3662 => x"04020101",
        3663 => x"05050505",
        3664 => x"05050202",
        3665 => x"02020202",
        3666 => x"05050505",
        3667 => x"06050505",
        3668 => x"05050206",
        3669 => x"03030202",
        3670 => x"02020206",
        3671 => x"02020202",
        3672 => x"02030502",
        3673 => x"06050505",
        3674 => x"05050206",
        3675 => x"02010304",
        3676 => x"04040404",
        3677 => x"04040404",
        3678 => x"04020103",
        3679 => x"02020202",
        3680 => x"02020202",
        3681 => x"02020202",
        3682 => x"02020202",
        3683 => x"02020202",
        3684 => x"02020202",
        3685 => x"02020202",
        3686 => x"02020202",
        3687 => x"02020202",
        3688 => x"02020202",
        3689 => x"02020202",
        3690 => x"02020202",
        3691 => x"02020202",
        3692 => x"02020202",
        3693 => x"02020202",
        3694 => x"02020202",
        3695 => x"02020202",
        3696 => x"02020202",
        3697 => x"02020202",
        3698 => x"02020202",
        3699 => x"02020202",
        3700 => x"02020202",
        3701 => x"02020202",
        3702 => x"02020202",
        3703 => x"02020202",
        3704 => x"02020202",
        3705 => x"02020202",
        3706 => x"02020202",
        3707 => x"02020202",
        3708 => x"02020202",
        3709 => x"02020202",
        3710 => x"02020202",

--			***** MAP *****

		
                --  MAP
        3711 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3712 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3713 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3714 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3715 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3716 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3717 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3718 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3719 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3720 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3721 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3722 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3723 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3724 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3725 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3726 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3727 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3728 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3729 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3730 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3731 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3732 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3733 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3734 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3735 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3736 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3737 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3738 => x"00000016", -- z: 0 rot: 0 ptr: 975
        3739 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3740 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3741 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3742 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3743 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3744 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3745 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3746 => x"00000038", -- z: 0 rot: 0 ptr: 1695
        3747 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3748 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3749 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3750 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3751 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3752 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3753 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3754 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3755 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3756 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3757 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3758 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3759 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3760 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3761 => x"00000038", -- z: 0 rot: 0 ptr: 1695
        3762 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3763 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3764 => x"00000003", -- z: 0 rot: 0 ptr: 471
        3765 => x"00000005", -- z: 0 rot: 0 ptr: 615
        3766 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3767 => x"00000003", -- z: 0 rot: 0 ptr: 471
        3768 => x"00000005", -- z: 0 rot: 0 ptr: 615
        3769 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3770 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3771 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3772 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3773 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3774 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3775 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3776 => x"00000038", -- z: 0 rot: 0 ptr: 1695
        3777 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3778 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3779 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3780 => x"00000015", -- z: 0 rot: 0 ptr: 903
        3781 => x"00000017", -- z: 0 rot: 0 ptr: 1047
        3782 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3783 => x"00000015", -- z: 0 rot: 0 ptr: 903
        3784 => x"00000017", -- z: 0 rot: 0 ptr: 1047
        3785 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3786 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3787 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3788 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3789 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3790 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3791 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3792 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3793 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3794 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3795 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3796 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3797 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3798 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3799 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3800 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3801 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3802 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3803 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3804 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3805 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3806 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3807 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3808 => x"00000026", -- z: 0 rot: 0 ptr: 1263
        3809 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3810 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3811 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3812 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3813 => x"00000003", -- z: 0 rot: 0 ptr: 471
        3814 => x"00000005", -- z: 0 rot: 0 ptr: 615
        3815 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3816 => x"00000003", -- z: 0 rot: 0 ptr: 471
        3817 => x"00000005", -- z: 0 rot: 0 ptr: 615
        3818 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3819 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3820 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3821 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3822 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3823 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3824 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3825 => x"00000026", -- z: 0 rot: 0 ptr: 1263
        3826 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3827 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3828 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3829 => x"00000015", -- z: 0 rot: 0 ptr: 903
        3830 => x"00000017", -- z: 0 rot: 0 ptr: 1047
        3831 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3832 => x"00000015", -- z: 0 rot: 0 ptr: 903
        3833 => x"00000017", -- z: 0 rot: 0 ptr: 1047
        3834 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3835 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3836 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3837 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3838 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3839 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3840 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3841 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3842 => x"00000026", -- z: 0 rot: 0 ptr: 1263
        3843 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3844 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3845 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3846 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3847 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3848 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3849 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3850 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3851 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3852 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3853 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3854 => x"00000002", -- z: 0 rot: 0 ptr: 399
        3855 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3856 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3857 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3858 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3859 => x"00000025", -- z: 0 rot: 0 ptr: 1191
        3860 => x"00000025", -- z: 0 rot: 0 ptr: 1191
        3861 => x"00000025", -- z: 0 rot: 0 ptr: 1191
        3862 => x"00000025", -- z: 0 rot: 0 ptr: 1191
        3863 => x"00000025", -- z: 0 rot: 0 ptr: 1191
        3864 => x"00000025", -- z: 0 rot: 0 ptr: 1191
        3865 => x"00000025", -- z: 0 rot: 0 ptr: 1191
        3866 => x"00000025", -- z: 0 rot: 0 ptr: 1191
        3867 => x"00000025", -- z: 0 rot: 0 ptr: 1191
        3868 => x"00000025", -- z: 0 rot: 0 ptr: 1191
        3869 => x"00000025", -- z: 0 rot: 0 ptr: 1191
        3870 => x"00000025", -- z: 0 rot: 0 ptr: 1191
        3871 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3872 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3873 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3874 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3875 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3876 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3877 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3878 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3879 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3880 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3881 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3882 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3883 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3884 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3885 => x"00000037", -- z: 0 rot: 0 ptr: 1623
        3886 => x"00000037", -- z: 0 rot: 0 ptr: 1623
		--stari je isao do 5438
		others => x"00000000"
	);


begin

	process(i_clk)
	begin
		if rising_edge(i_clk) then
			-- memory write --
			if i_we = '1' then
				mem(to_integer(unsigned(i_w_addr))) <= i_data;
			end if;
			-- memory read -- 
			o_data <= mem(to_integer(unsigned(i_r_addr)));
			
		end if; 
	end process;

end architecture arch;