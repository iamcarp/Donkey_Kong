
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity ram is
	generic
	(
		DATA_WIDTH : natural := 32;		    -- 4 byte one line of memory
		ADDR_WIDTH : natural := 13			    -- 24576 bytes size of memory
	);

	port(
		i_clk    : in  std_logic;
		i_r_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		i_data   : in  std_logic_vector(DATA_WIDTH-1 downto 0);
		i_we     : in  std_logic;
		i_w_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		o_data   : out std_logic_vector(DATA_WIDTH-1 downto 0)
	);
end entity ram;

architecture arch of ram is

	type ram_t is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(DATA_WIDTH-1 downto 0);


-- GENERATED BY BC_MEM_PACKER

-- DATE: Thu May 18 16:01:02 2017

	signal mem : ram_t := (

--			***** COLOR PALLETE *****

		-- fellas
		0 =>	x"000C4CC8",
		1 =>	x"00A8D8FC",
		2 =>	x"00000000",
		3 =>	x"00EC3820",
		4 =>	x"0000A800",
		5 =>	x"00FCFCFC",
		6 =>	x"00747474",
		7 =>	x"00C0C0C0",
--      Link colors
        8 =>    x"00303030",
        9 =>    x"000CCB83",
        10 =>   x"002C98D8",
        11 =>   x"00004B7B",
        12 =>   x"00FFD9D9",
        13 =>   x"00003299",
        14 =>   x"00B1DFF8",
        15 =>   x"00FFFFFF",
        16 =>   x"008E0018",
        17 =>   x"00FF898E",
        18 =>   x"00000000",
        19 =>   x"00006E8A",
        20 =>   x"00002E55",
        21 =>   x"00CBC74D",
        22 =>   x"00E32F47",
        23 =>   x"00173B00",
        24 =>   x"00007A3E",
        25 =>   x"007ED14A",
        26 =>   x"0000311D",
        27 =>   x"0000675B",
        28 =>   x"000AB4B9",
        29 =>   x"00003D00",
        30 =>   x"00008200",
        31 =>   x"003FD65B",
        32 =>   x"00656565",
        33 =>   x"00B9B9B9",
        34 =>   x"00AFAFAF",
-- 		enemie colors
		35 =>	x"00c0c0c0",
		36 => 	x"000038f8",
		37 => 	x"00bc0000",
		38 =>	x"00ff8868",
		39 => 	x"00ffffff",
																															-- map colors

																															40=> x"00000000",
																															41=> x"00bc0000",
																															42=> x"00d8e800",
																															43=> x"00010100",
																															44=> x"00010000",
																															45=> x"0044a0fc",

							46 => x"00523900",
							47 => x"00271900",
							48 => x"00080400",
							49 => x"00010000",
							50 => x"00d8e800",
							51 => x"00000a00",
							52 => x"0000d600",
							53 => x"00020202",
							54 => x"00010101",
							55 => x"00010100",
							56 => x"00030600",
							57 => x"00105ce4",
							58 => x"0044a0fc",
							59 => x"00bc0000",
							60 => x"005800e4",
							61 => x"00020100",
							62 => x"00f85800",
		63 =>	x"003199FF", -- Unused

            --  ADDED SPRITES HERE
          -- RUPEE SPRITE
		64 => x"0202020F",
		65 => x"3C020202",
		66 => x"02020202",
		67 => x"02020202",
		68 => x"02020F0F",
		69 => x"3C3C0202",
		70 => x"02020202",
		71 => x"02020202",
		72 => x"020F0F0F",
		73 => x"3C3C3C02",
		74 => x"02020202",
		75 => x"02020202",
		76 => x"0F3C0F3C",
		77 => x"023C023C",
		78 => x"02020202",
		79 => x"02020202",
		80 => x"0F0F3C3C",
		81 => x"3C023C3C",
		82 => x"02020202",
		83 => x"02020202",
		84 => x"0F0F3C3C",
		85 => x"3C023C3C",
		86 => x"02020202",
		87 => x"02020202",
		88 => x"0F0F3C3C",
		89 => x"3C023C3C",
		90 => x"02020202",
		91 => x"02020202",
		92 => x"0F0F3C3C",
		93 => x"3C023C3C",
		94 => x"02020202",
		95 => x"02020202",
		96 => x"0F0F3C3C",
		97 => x"3C023C3C",
		98 => x"02020202",
		99 => x"02020202",
		100 => x"0F0F3C3C",
		101 => x"3C023C3C",
		102 => x"02020202",
		103 => x"02020202",
		104 => x"0F0F3C3C",
		105 => x"3C023C3C",
		106 => x"02020202",
		107 => x"02020202",
		108 => x"0F3C0F3C",
		109 => x"3C023C3C",
		110 => x"02020202",
		111 => x"02020202",
		112 => x"3C3C3C0F",
		113 => x"023C023C",
		114 => x"02020202",
		115 => x"02020202",
		116 => x"023C3C3C",
		117 => x"3C3C3C02",
		118 => x"02020202",
		119 => x"02020202",
		120 => x"02023C3C",
		121 => x"3C3C0202",
		122 => x"02020202",
		123 => x"02020202",
		124 => x"0202023C",
		125 => x"3C020202",
		126 => x"02020202",
		127 => x"02020202",

          -- BOMB SPRITE
		128 => x"02020202",
		129 => x"020F0202",
		130 => x"02020202",
		131 => x"02020202",
		132 => x"02020202",
		133 => x"020F0202",
		134 => x"02020202",
		135 => x"02020202",
		136 => x"02020202",
		137 => x"02020F02",
		138 => x"02020202",
		139 => x"02020202",
		140 => x"02020202",
		141 => x"0202020F",
		142 => x"02020202",
		143 => x"02020202",
		144 => x"02020202",
		145 => x"0202020F",
		146 => x"02020202",
		147 => x"02020202",
		148 => x"02020202",
		149 => x"02020F02",
		150 => x"02020202",
		151 => x"02020202",
		152 => x"02020D0D",
		153 => x"0D0D0202",
		154 => x"02020202",
		155 => x"02020202",
		156 => x"020D2E2E",
		157 => x"0D0D0D02",
		158 => x"02020202",
		159 => x"02020202",
		160 => x"0D2E0F2E",
		161 => x"0D0D0D0D",
		162 => x"02020202",
		163 => x"02020202",
		164 => x"0D2E2E0D",
		165 => x"0D0D0D0D",
		166 => x"02020202",
		167 => x"02020202",
		168 => x"0D0D0D0D",
		169 => x"0D0D0D0D",
		170 => x"02020202",
		171 => x"02020202",
		172 => x"0D0D0D0D",
		173 => x"0D0D0D0D",
		174 => x"02020202",
		175 => x"02020202",
		176 => x"020D0D0D",
		177 => x"0D0D0D02",
		178 => x"02020202",
		179 => x"02020202",
		180 => x"02020D0D",
		181 => x"0D0D0202",
		182 => x"02020202",
		183 => x"02020202",
		184 => x"02020202",
		185 => x"02020202",
		186 => x"02020202",
		187 => x"02020202",
		188 => x"02020202",
		189 => x"02020202",
		190 => x"02020202",
		191 => x"02020202",

--			***** 16x16 IMAGES *****
--			OVERWORLD SPRITES


						--  sprite 0
		255 => x"00000000",		-- colors: 40, 40, 40, 40
		256 => x"00000000",		-- colors: 40, 40, 40, 40
		257 => x"00000000",		-- colors: 40, 40, 40, 40
		258 => x"00000000",		-- colors: 40, 40, 40, 40
		259 => x"29292929",		-- colors: 41, 41, 41, 41
		260 => x"29292929",		-- colors: 41, 41, 41, 41
		261 => x"29292929",		-- colors: 41, 41, 41, 41
		262 => x"29292929",		-- colors: 41, 41, 41, 41
		263 => x"00002A2A",		-- colors: 40, 40, 42, 42
		264 => x"2A2A0000",		-- colors: 42, 42, 40, 40
		265 => x"00002A2A",		-- colors: 40, 40, 42, 42
		266 => x"2A2A0000",		-- colors: 42, 42, 40, 40
		267 => x"002A2A2A",		-- colors: 40, 42, 42, 42
		268 => x"2A2A2A00",		-- colors: 42, 42, 42, 40
		269 => x"002A2A2A",		-- colors: 40, 42, 42, 42
		270 => x"2A2A2A00",		-- colors: 42, 42, 42, 40
		271 => x"002A2A2A",		-- colors: 40, 42, 42, 42
		272 => x"2A2A2A00",		-- colors: 42, 42, 42, 40
		273 => x"002A2A2A",		-- colors: 40, 42, 42, 42
		274 => x"2A2A2A00",		-- colors: 42, 42, 42, 40
		275 => x"00002A2A",		-- colors: 40, 40, 42, 42
		276 => x"2A2A0000",		-- colors: 42, 42, 40, 40
		277 => x"00002A2A",		-- colors: 40, 40, 42, 42
		278 => x"2A2A0000",		-- colors: 42, 42, 40, 40
		279 => x"00000000",		-- colors: 40, 40, 40, 40
		280 => x"00000000",		-- colors: 40, 40, 40, 40
		281 => x"00000000",		-- colors: 40, 40, 40, 40
		282 => x"00000000",		-- colors: 40, 40, 40, 40
		283 => x"29292929",		-- colors: 41, 41, 41, 41
		284 => x"29292929",		-- colors: 41, 41, 41, 41
		285 => x"29292929",		-- colors: 41, 41, 41, 41
		286 => x"29292929",		-- colors: 41, 41, 41, 41
		287 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		288 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		289 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		290 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		291 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		292 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		293 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		294 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		295 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		296 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		297 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		298 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		299 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		300 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		301 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		302 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		303 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		304 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		305 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		306 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		307 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		308 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		309 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		310 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		311 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		312 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		313 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		314 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		315 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		316 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		317 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		318 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42

						--  sprite 1
		319 => x"00000000",		-- colors: 40, 40, 40, 40
		320 => x"00000000",		-- colors: 40, 40, 40, 40
		321 => x"00000000",		-- colors: 40, 40, 40, 40
		322 => x"00000000",		-- colors: 40, 40, 40, 40
		323 => x"00000000",		-- colors: 40, 40, 40, 40
		324 => x"00000000",		-- colors: 40, 40, 40, 40
		325 => x"00000000",		-- colors: 40, 40, 40, 40
		326 => x"00000000",		-- colors: 40, 40, 40, 40
		327 => x"00000000",		-- colors: 40, 40, 40, 40
		328 => x"00000000",		-- colors: 40, 40, 40, 40
		329 => x"00000000",		-- colors: 40, 40, 40, 40
		330 => x"00000000",		-- colors: 40, 40, 40, 40
		331 => x"00000000",		-- colors: 40, 40, 40, 40
		332 => x"00000000",		-- colors: 40, 40, 40, 40
		333 => x"00000000",		-- colors: 40, 40, 40, 40
		334 => x"00000000",		-- colors: 40, 40, 40, 40
		335 => x"00000000",		-- colors: 40, 40, 40, 40
		336 => x"00000000",		-- colors: 40, 40, 40, 40
		337 => x"00000000",		-- colors: 40, 40, 40, 40
		338 => x"00000000",		-- colors: 40, 40, 40, 40
		339 => x"00000000",		-- colors: 40, 40, 40, 40
		340 => x"00000000",		-- colors: 40, 40, 40, 40
		341 => x"00000000",		-- colors: 40, 40, 40, 40
		342 => x"00000000",		-- colors: 40, 40, 40, 40
		343 => x"00000000",		-- colors: 40, 40, 40, 40
		344 => x"00000000",		-- colors: 40, 40, 40, 40
		345 => x"00000000",		-- colors: 40, 40, 40, 40
		346 => x"00000000",		-- colors: 40, 40, 40, 40
		347 => x"00000000",		-- colors: 40, 40, 40, 40
		348 => x"00000000",		-- colors: 40, 40, 40, 40
		349 => x"00000000",		-- colors: 40, 40, 40, 40
		350 => x"00000000",		-- colors: 40, 40, 40, 40
		351 => x"29292929",		-- colors: 41, 41, 41, 41
		352 => x"29292929",		-- colors: 41, 41, 41, 41
		353 => x"29292929",		-- colors: 41, 41, 41, 41
		354 => x"29292929",		-- colors: 41, 41, 41, 41
		355 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		356 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		357 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		358 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		359 => x"29290000",		-- colors: 41, 41, 40, 40
		360 => x"00002929",		-- colors: 40, 40, 41, 41
		361 => x"29290000",		-- colors: 41, 41, 40, 40
		362 => x"00002929",		-- colors: 40, 40, 41, 41
		363 => x"29000000",		-- colors: 41, 40, 40, 40
		364 => x"00000029",		-- colors: 40, 40, 40, 41
		365 => x"29000000",		-- colors: 41, 40, 40, 40
		366 => x"00000029",		-- colors: 40, 40, 40, 41
		367 => x"29000000",		-- colors: 41, 40, 40, 40
		368 => x"00000029",		-- colors: 40, 40, 40, 41
		369 => x"29000000",		-- colors: 41, 40, 40, 40
		370 => x"00000029",		-- colors: 40, 40, 40, 41
		371 => x"29290000",		-- colors: 41, 41, 40, 40
		372 => x"00002929",		-- colors: 40, 40, 41, 41
		373 => x"29290000",		-- colors: 41, 41, 40, 40
		374 => x"00002929",		-- colors: 40, 40, 41, 41
		375 => x"29292929",		-- colors: 41, 41, 41, 41
		376 => x"29292929",		-- colors: 41, 41, 41, 41
		377 => x"29292929",		-- colors: 41, 41, 41, 41
		378 => x"29292929",		-- colors: 41, 41, 41, 41
		379 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		380 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		381 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		382 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42

						--  sprite 2
		383 => x"00000000",		-- colors: 40, 40, 40, 40
		384 => x"00000000",		-- colors: 40, 40, 40, 40
		385 => x"29000000",		-- colors: 41, 40, 40, 40
		386 => x"00000029",		-- colors: 40, 40, 40, 41
		387 => x"00000000",		-- colors: 40, 40, 40, 40
		388 => x"00000000",		-- colors: 40, 40, 40, 40
		389 => x"29292929",		-- colors: 41, 41, 41, 41
		390 => x"29292929",		-- colors: 41, 41, 41, 41
		391 => x"00000000",		-- colors: 40, 40, 40, 40
		392 => x"00000000",		-- colors: 40, 40, 40, 40
		393 => x"29000000",		-- colors: 41, 40, 40, 40
		394 => x"00000029",		-- colors: 40, 40, 40, 41
		395 => x"00000000",		-- colors: 40, 40, 40, 40
		396 => x"00000000",		-- colors: 40, 40, 40, 40
		397 => x"29000000",		-- colors: 41, 40, 40, 40
		398 => x"00000029",		-- colors: 40, 40, 40, 41
		399 => x"00000000",		-- colors: 40, 40, 40, 40
		400 => x"00000000",		-- colors: 40, 40, 40, 40
		401 => x"29000000",		-- colors: 41, 40, 40, 40
		402 => x"00000029",		-- colors: 40, 40, 40, 41
		403 => x"00000000",		-- colors: 40, 40, 40, 40
		404 => x"00000000",		-- colors: 40, 40, 40, 40
		405 => x"29292929",		-- colors: 41, 41, 41, 41
		406 => x"29292929",		-- colors: 41, 41, 41, 41
		407 => x"00000000",		-- colors: 40, 40, 40, 40
		408 => x"00000000",		-- colors: 40, 40, 40, 40
		409 => x"29000000",		-- colors: 41, 40, 40, 40
		410 => x"00000029",		-- colors: 40, 40, 40, 41
		411 => x"00000000",		-- colors: 40, 40, 40, 40
		412 => x"00000000",		-- colors: 40, 40, 40, 40
		413 => x"29000000",		-- colors: 41, 40, 40, 40
		414 => x"00000029",		-- colors: 40, 40, 40, 41
		415 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		416 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		417 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		418 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		419 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
		420 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
		421 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
		422 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
		423 => x"2A2A0000",		-- colors: 42, 42, 40, 40
		424 => x"00002A2A",		-- colors: 40, 40, 42, 42
		425 => x"2A2A0000",		-- colors: 42, 42, 40, 40
		426 => x"00002A2A",		-- colors: 40, 40, 42, 42
		427 => x"2A000000",		-- colors: 42, 40, 40, 40
		428 => x"0000002A",		-- colors: 40, 40, 40, 42
		429 => x"2A000000",		-- colors: 42, 40, 40, 40
		430 => x"0000002A",		-- colors: 40, 40, 40, 42
		431 => x"2A000000",		-- colors: 42, 40, 40, 40
		432 => x"0000002A",		-- colors: 40, 40, 40, 42
		433 => x"2A000000",		-- colors: 42, 40, 40, 40
		434 => x"0000002A",		-- colors: 40, 40, 40, 42
		435 => x"2A2A0000",		-- colors: 42, 42, 40, 40
		436 => x"00002A2A",		-- colors: 40, 40, 42, 42
		437 => x"2A2A0000",		-- colors: 42, 42, 40, 40
		438 => x"00002A2A",		-- colors: 40, 40, 42, 42
		439 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		440 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		441 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		442 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		443 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
		444 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
		445 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
		446 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43

						--  sprite 3
		447 => x"00292929",		-- colors: 40, 41, 41, 41
		448 => x"29292900",		-- colors: 41, 41, 41, 40
		449 => x"29292929",		-- colors: 41, 41, 41, 41
		450 => x"29292929",		-- colors: 41, 41, 41, 41
		451 => x"00000000",		-- colors: 40, 40, 40, 40
		452 => x"00000000",		-- colors: 40, 40, 40, 40
		453 => x"29292929",		-- colors: 41, 41, 41, 41
		454 => x"29292929",		-- colors: 41, 41, 41, 41
		455 => x"00292929",		-- colors: 40, 41, 41, 41
		456 => x"29292900",		-- colors: 41, 41, 41, 40
		457 => x"29292929",		-- colors: 41, 41, 41, 41
		458 => x"29292929",		-- colors: 41, 41, 41, 41
		459 => x"00292929",		-- colors: 40, 41, 41, 41
		460 => x"29292900",		-- colors: 41, 41, 41, 40
		461 => x"29292929",		-- colors: 41, 41, 41, 41
		462 => x"29292929",		-- colors: 41, 41, 41, 41
		463 => x"00292929",		-- colors: 40, 41, 41, 41
		464 => x"29292900",		-- colors: 41, 41, 41, 40
		465 => x"29292929",		-- colors: 41, 41, 41, 41
		466 => x"29292929",		-- colors: 41, 41, 41, 41
		467 => x"00000000",		-- colors: 40, 40, 40, 40
		468 => x"00000000",		-- colors: 40, 40, 40, 40
		469 => x"29292929",		-- colors: 41, 41, 41, 41
		470 => x"29292929",		-- colors: 41, 41, 41, 41
		471 => x"00292929",		-- colors: 40, 41, 41, 41
		472 => x"29292900",		-- colors: 41, 41, 41, 40
		473 => x"29292929",		-- colors: 41, 41, 41, 41
		474 => x"29292929",		-- colors: 41, 41, 41, 41
		475 => x"00292929",		-- colors: 40, 41, 41, 41
		476 => x"29292900",		-- colors: 41, 41, 41, 40
		477 => x"29292929",		-- colors: 41, 41, 41, 41
		478 => x"29292929",		-- colors: 41, 41, 41, 41
		479 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		480 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		481 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		482 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		483 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
		484 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
		485 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
		486 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
		487 => x"2A2A2929",		-- colors: 42, 42, 41, 41
		488 => x"29292A2A",		-- colors: 41, 41, 42, 42
		489 => x"2A2A2929",		-- colors: 42, 42, 41, 41
		490 => x"29292A2A",		-- colors: 41, 41, 42, 42
		491 => x"2A292929",		-- colors: 42, 41, 41, 41
		492 => x"2929292A",		-- colors: 41, 41, 41, 42
		493 => x"2A292929",		-- colors: 42, 41, 41, 41
		494 => x"2929292A",		-- colors: 41, 41, 41, 42
		495 => x"2A292929",		-- colors: 42, 41, 41, 41
		496 => x"2929292A",		-- colors: 41, 41, 41, 42
		497 => x"2A292929",		-- colors: 42, 41, 41, 41
		498 => x"2929292A",		-- colors: 41, 41, 41, 42
		499 => x"2A2A2929",		-- colors: 42, 42, 41, 41
		500 => x"29292A2A",		-- colors: 41, 41, 42, 42
		501 => x"2A2A2929",		-- colors: 42, 42, 41, 41
		502 => x"29292A2A",		-- colors: 41, 41, 42, 42
		503 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		504 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		505 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		506 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		507 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
		508 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
		509 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
		510 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43

						--  sprite 4
		511 => x"00292929",		-- colors: 40, 41, 41, 41
		512 => x"29292900",		-- colors: 41, 41, 41, 40
		513 => x"29292929",		-- colors: 41, 41, 41, 41
		514 => x"29292929",		-- colors: 41, 41, 41, 41
		515 => x"00000000",		-- colors: 40, 40, 40, 40
		516 => x"00000000",		-- colors: 40, 40, 40, 40
		517 => x"29292929",		-- colors: 41, 41, 41, 41
		518 => x"29292929",		-- colors: 41, 41, 41, 41
		519 => x"00292929",		-- colors: 40, 41, 41, 41
		520 => x"29292900",		-- colors: 41, 41, 41, 40
		521 => x"29292929",		-- colors: 41, 41, 41, 41
		522 => x"29292929",		-- colors: 41, 41, 41, 41
		523 => x"00292929",		-- colors: 40, 41, 41, 41
		524 => x"29292900",		-- colors: 41, 41, 41, 40
		525 => x"29292929",		-- colors: 41, 41, 41, 41
		526 => x"29292929",		-- colors: 41, 41, 41, 41
		527 => x"00292929",		-- colors: 40, 41, 41, 41
		528 => x"29292900",		-- colors: 41, 41, 41, 40
		529 => x"29292929",		-- colors: 41, 41, 41, 41
		530 => x"29292929",		-- colors: 41, 41, 41, 41
		531 => x"00000000",		-- colors: 40, 40, 40, 40
		532 => x"00000000",		-- colors: 40, 40, 40, 40
		533 => x"29292929",		-- colors: 41, 41, 41, 41
		534 => x"29292929",		-- colors: 41, 41, 41, 41
		535 => x"00292929",		-- colors: 40, 41, 41, 41
		536 => x"29292900",		-- colors: 41, 41, 41, 40
		537 => x"29292929",		-- colors: 41, 41, 41, 41
		538 => x"29292929",		-- colors: 41, 41, 41, 41
		539 => x"00292929",		-- colors: 40, 41, 41, 41
		540 => x"29292900",		-- colors: 41, 41, 41, 40
		541 => x"29292929",		-- colors: 41, 41, 41, 41
		542 => x"29292929",		-- colors: 41, 41, 41, 41
		543 => x"00292929",		-- colors: 40, 41, 41, 41
		544 => x"29292900",		-- colors: 41, 41, 41, 40
		545 => x"29292929",		-- colors: 41, 41, 41, 41
		546 => x"29292929",		-- colors: 41, 41, 41, 41
		547 => x"00000000",		-- colors: 40, 40, 40, 40
		548 => x"00000000",		-- colors: 40, 40, 40, 40
		549 => x"29292929",		-- colors: 41, 41, 41, 41
		550 => x"29292929",		-- colors: 41, 41, 41, 41
		551 => x"00292929",		-- colors: 40, 41, 41, 41
		552 => x"29292900",		-- colors: 41, 41, 41, 40
		553 => x"29292929",		-- colors: 41, 41, 41, 41
		554 => x"29292929",		-- colors: 41, 41, 41, 41
		555 => x"00292929",		-- colors: 40, 41, 41, 41
		556 => x"29292900",		-- colors: 41, 41, 41, 40
		557 => x"29292929",		-- colors: 41, 41, 41, 41
		558 => x"29292929",		-- colors: 41, 41, 41, 41
		559 => x"00292929",		-- colors: 40, 41, 41, 41
		560 => x"29292900",		-- colors: 41, 41, 41, 40
		561 => x"29292929",		-- colors: 41, 41, 41, 41
		562 => x"29292929",		-- colors: 41, 41, 41, 41
		563 => x"00000000",		-- colors: 40, 40, 40, 40
		564 => x"00000000",		-- colors: 40, 40, 40, 40
		565 => x"29292929",		-- colors: 41, 41, 41, 41
		566 => x"29292929",		-- colors: 41, 41, 41, 41
		567 => x"00292929",		-- colors: 40, 41, 41, 41
		568 => x"29292900",		-- colors: 41, 41, 41, 40
		569 => x"29292929",		-- colors: 41, 41, 41, 41
		570 => x"29292929",		-- colors: 41, 41, 41, 41
		571 => x"00292929",		-- colors: 40, 41, 41, 41
		572 => x"29292900",		-- colors: 41, 41, 41, 40
		573 => x"29292929",		-- colors: 41, 41, 41, 41
		574 => x"29292929",		-- colors: 41, 41, 41, 41

						--  sprite 5
		575 => x"00000000",		-- colors: 40, 40, 40, 40
		576 => x"00000000",		-- colors: 40, 40, 40, 40
		577 => x"29000000",		-- colors: 41, 40, 40, 40
		578 => x"00000029",		-- colors: 40, 40, 40, 41
		579 => x"00000000",		-- colors: 40, 40, 40, 40
		580 => x"00000000",		-- colors: 40, 40, 40, 40
		581 => x"29292929",		-- colors: 41, 41, 41, 41
		582 => x"29292929",		-- colors: 41, 41, 41, 41
		583 => x"00000000",		-- colors: 40, 40, 40, 40
		584 => x"00000000",		-- colors: 40, 40, 40, 40
		585 => x"29000000",		-- colors: 41, 40, 40, 40
		586 => x"00000029",		-- colors: 40, 40, 40, 41
		587 => x"00000000",		-- colors: 40, 40, 40, 40
		588 => x"00000000",		-- colors: 40, 40, 40, 40
		589 => x"29000000",		-- colors: 41, 40, 40, 40
		590 => x"00000029",		-- colors: 40, 40, 40, 41
		591 => x"00000000",		-- colors: 40, 40, 40, 40
		592 => x"00000000",		-- colors: 40, 40, 40, 40
		593 => x"29000000",		-- colors: 41, 40, 40, 40
		594 => x"00000029",		-- colors: 40, 40, 40, 41
		595 => x"00000000",		-- colors: 40, 40, 40, 40
		596 => x"00000000",		-- colors: 40, 40, 40, 40
		597 => x"29292929",		-- colors: 41, 41, 41, 41
		598 => x"29292929",		-- colors: 41, 41, 41, 41
		599 => x"00000000",		-- colors: 40, 40, 40, 40
		600 => x"00000000",		-- colors: 40, 40, 40, 40
		601 => x"29000000",		-- colors: 41, 40, 40, 40
		602 => x"00000029",		-- colors: 40, 40, 40, 41
		603 => x"00000000",		-- colors: 40, 40, 40, 40
		604 => x"00000000",		-- colors: 40, 40, 40, 40
		605 => x"29000000",		-- colors: 41, 40, 40, 40
		606 => x"00000029",		-- colors: 40, 40, 40, 41
		607 => x"00000000",		-- colors: 40, 40, 40, 40
		608 => x"00000000",		-- colors: 40, 40, 40, 40
		609 => x"29000000",		-- colors: 41, 40, 40, 40
		610 => x"00000029",		-- colors: 40, 40, 40, 41
		611 => x"00000000",		-- colors: 40, 40, 40, 40
		612 => x"00000000",		-- colors: 40, 40, 40, 40
		613 => x"29292929",		-- colors: 41, 41, 41, 41
		614 => x"29292929",		-- colors: 41, 41, 41, 41
		615 => x"00000000",		-- colors: 40, 40, 40, 40
		616 => x"00000000",		-- colors: 40, 40, 40, 40
		617 => x"29000000",		-- colors: 41, 40, 40, 40
		618 => x"00000029",		-- colors: 40, 40, 40, 41
		619 => x"00000000",		-- colors: 40, 40, 40, 40
		620 => x"00000000",		-- colors: 40, 40, 40, 40
		621 => x"29000000",		-- colors: 41, 40, 40, 40
		622 => x"00000029",		-- colors: 40, 40, 40, 41
		623 => x"00000000",		-- colors: 40, 40, 40, 40
		624 => x"00000000",		-- colors: 40, 40, 40, 40
		625 => x"29000000",		-- colors: 41, 40, 40, 40
		626 => x"00000029",		-- colors: 40, 40, 40, 41
		627 => x"00000000",		-- colors: 40, 40, 40, 40
		628 => x"00000000",		-- colors: 40, 40, 40, 40
		629 => x"29292929",		-- colors: 41, 41, 41, 41
		630 => x"29292929",		-- colors: 41, 41, 41, 41
		631 => x"00000000",		-- colors: 40, 40, 40, 40
		632 => x"00000000",		-- colors: 40, 40, 40, 40
		633 => x"29000000",		-- colors: 41, 40, 40, 40
		634 => x"00000029",		-- colors: 40, 40, 40, 41
		635 => x"00000000",		-- colors: 40, 40, 40, 40
		636 => x"00000000",		-- colors: 40, 40, 40, 40
		637 => x"29000000",		-- colors: 41, 40, 40, 40
		638 => x"00000029",		-- colors: 40, 40, 40, 41

						--  sprite 6
		639 => x"00000000",		-- colors: 40, 40, 40, 40
		640 => x"00000000",		-- colors: 40, 40, 40, 40
		641 => x"00000000",		-- colors: 40, 40, 40, 40
		642 => x"00000000",		-- colors: 40, 40, 40, 40
		643 => x"00000000",		-- colors: 40, 40, 40, 40
		644 => x"00000000",		-- colors: 40, 40, 40, 40
		645 => x"00000000",		-- colors: 40, 40, 40, 40
		646 => x"00000000",		-- colors: 40, 40, 40, 40
		647 => x"00000000",		-- colors: 40, 40, 40, 40
		648 => x"00000000",		-- colors: 40, 40, 40, 40
		649 => x"00000000",		-- colors: 40, 40, 40, 40
		650 => x"00000000",		-- colors: 40, 40, 40, 40
		651 => x"00000000",		-- colors: 40, 40, 40, 40
		652 => x"00000000",		-- colors: 40, 40, 40, 40
		653 => x"00000000",		-- colors: 40, 40, 40, 40
		654 => x"00000000",		-- colors: 40, 40, 40, 40
		655 => x"00000000",		-- colors: 40, 40, 40, 40
		656 => x"00000000",		-- colors: 40, 40, 40, 40
		657 => x"00000000",		-- colors: 40, 40, 40, 40
		658 => x"00000000",		-- colors: 40, 40, 40, 40
		659 => x"00000000",		-- colors: 40, 40, 40, 40
		660 => x"00000000",		-- colors: 40, 40, 40, 40
		661 => x"00000000",		-- colors: 40, 40, 40, 40
		662 => x"00000000",		-- colors: 40, 40, 40, 40
		663 => x"00000000",		-- colors: 40, 40, 40, 40
		664 => x"00000000",		-- colors: 40, 40, 40, 40
		665 => x"00000000",		-- colors: 40, 40, 40, 40
		666 => x"00000000",		-- colors: 40, 40, 40, 40
		667 => x"00000000",		-- colors: 40, 40, 40, 40
		668 => x"00000000",		-- colors: 40, 40, 40, 40
		669 => x"00000000",		-- colors: 40, 40, 40, 40
		670 => x"00000000",		-- colors: 40, 40, 40, 40
		671 => x"00000000",		-- colors: 40, 40, 40, 40
		672 => x"00000000",		-- colors: 40, 40, 40, 40
		673 => x"00000000",		-- colors: 40, 40, 40, 40
		674 => x"00000000",		-- colors: 40, 40, 40, 40
		675 => x"00000000",		-- colors: 40, 40, 40, 40
		676 => x"00000000",		-- colors: 40, 40, 40, 40
		677 => x"00000000",		-- colors: 40, 40, 40, 40
		678 => x"00000000",		-- colors: 40, 40, 40, 40
		679 => x"00000000",		-- colors: 40, 40, 40, 40
		680 => x"00000000",		-- colors: 40, 40, 40, 40
		681 => x"00000000",		-- colors: 40, 40, 40, 40
		682 => x"00000000",		-- colors: 40, 40, 40, 40
		683 => x"00000000",		-- colors: 40, 40, 40, 40
		684 => x"00000000",		-- colors: 40, 40, 40, 40
		685 => x"00000000",		-- colors: 40, 40, 40, 40
		686 => x"00000000",		-- colors: 40, 40, 40, 40
		687 => x"00000000",		-- colors: 40, 40, 40, 40
		688 => x"00000000",		-- colors: 40, 40, 40, 40
		689 => x"00000000",		-- colors: 40, 40, 40, 40
		690 => x"00000000",		-- colors: 40, 40, 40, 40
		691 => x"00000000",		-- colors: 40, 40, 40, 40
		692 => x"00000000",		-- colors: 40, 40, 40, 40
		693 => x"00000000",		-- colors: 40, 40, 40, 40
		694 => x"00000000",		-- colors: 40, 40, 40, 40
		695 => x"00000000",		-- colors: 40, 40, 40, 40
		696 => x"00000000",		-- colors: 40, 40, 40, 40
		697 => x"00000000",		-- colors: 40, 40, 40, 40
		698 => x"00000000",		-- colors: 40, 40, 40, 40
		699 => x"00000000",		-- colors: 40, 40, 40, 40
		700 => x"00000000",		-- colors: 40, 40, 40, 40
		701 => x"00000000",		-- colors: 40, 40, 40, 40
		702 => x"00000000",		-- colors: 40, 40, 40, 40

						--  sprite 7
		703 => x"00000000",		-- colors: 40, 40, 40, 40
		704 => x"00000000",		-- colors: 40, 40, 40, 40
		705 => x"00000000",		-- colors: 40, 40, 40, 40
		706 => x"00000000",		-- colors: 40, 40, 40, 40
		707 => x"29292929",		-- colors: 41, 41, 41, 41
		708 => x"29292929",		-- colors: 41, 41, 41, 41
		709 => x"29292929",		-- colors: 41, 41, 41, 41
		710 => x"29292929",		-- colors: 41, 41, 41, 41
		711 => x"00002A2A",		-- colors: 40, 40, 42, 42
		712 => x"2A2A0000",		-- colors: 42, 42, 40, 40
		713 => x"00002A2A",		-- colors: 40, 40, 42, 42
		714 => x"2A2A0000",		-- colors: 42, 42, 40, 40
		715 => x"002A2A2A",		-- colors: 40, 42, 42, 42
		716 => x"2A2A2A00",		-- colors: 42, 42, 42, 40
		717 => x"002A2A2A",		-- colors: 40, 42, 42, 42
		718 => x"2A2A2A00",		-- colors: 42, 42, 42, 40
		719 => x"002A2A2A",		-- colors: 40, 42, 42, 42
		720 => x"2A2A2A00",		-- colors: 42, 42, 42, 40
		721 => x"002A2A2A",		-- colors: 40, 42, 42, 42
		722 => x"2A2A2A00",		-- colors: 42, 42, 42, 40
		723 => x"00002A2A",		-- colors: 40, 40, 42, 42
		724 => x"2A2A0000",		-- colors: 42, 42, 40, 40
		725 => x"00002A2A",		-- colors: 40, 40, 42, 42
		726 => x"2A2A0000",		-- colors: 42, 42, 40, 40
		727 => x"00000000",		-- colors: 40, 40, 40, 40
		728 => x"00000000",		-- colors: 40, 40, 40, 40
		729 => x"00000000",		-- colors: 40, 40, 40, 40
		730 => x"00000000",		-- colors: 40, 40, 40, 40
		731 => x"29292929",		-- colors: 41, 41, 41, 41
		732 => x"29292929",		-- colors: 41, 41, 41, 41
		733 => x"29292929",		-- colors: 41, 41, 41, 41
		734 => x"29292929",		-- colors: 41, 41, 41, 41
		735 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		736 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		737 => x"2B2A2A2A",		-- colors: 43, 42, 42, 42
		738 => x"2A2A2A2B",		-- colors: 42, 42, 42, 43
		739 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		740 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		741 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
		742 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
		743 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		744 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		745 => x"2B2A2A2A",		-- colors: 43, 42, 42, 42
		746 => x"2A2A2A2B",		-- colors: 42, 42, 42, 43
		747 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		748 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		749 => x"2B2A2A2A",		-- colors: 43, 42, 42, 42
		750 => x"2A2A2A2B",		-- colors: 42, 42, 42, 43
		751 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		752 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		753 => x"2B2A2A2A",		-- colors: 43, 42, 42, 42
		754 => x"2A2A2A2B",		-- colors: 42, 42, 42, 43
		755 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		756 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		757 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
		758 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
		759 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		760 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		761 => x"2B2A2A2A",		-- colors: 43, 42, 42, 42
		762 => x"2A2A2A2B",		-- colors: 42, 42, 42, 43
		763 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		764 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		765 => x"2B2A2A2A",		-- colors: 43, 42, 42, 42
		766 => x"2A2A2A2B",		-- colors: 42, 42, 42, 43

						--  sprite 8
		767 => x"00000000",		-- colors: 40, 40, 40, 40
		768 => x"00000000",		-- colors: 40, 40, 40, 40
		769 => x"00000000",		-- colors: 40, 40, 40, 40
		770 => x"00000000",		-- colors: 40, 40, 40, 40
		771 => x"29292929",		-- colors: 41, 41, 41, 41
		772 => x"29292929",		-- colors: 41, 41, 41, 41
		773 => x"29292929",		-- colors: 41, 41, 41, 41
		774 => x"29292929",		-- colors: 41, 41, 41, 41
		775 => x"00002A2A",		-- colors: 40, 40, 42, 42
		776 => x"2A2A0000",		-- colors: 42, 42, 40, 40
		777 => x"00002A2A",		-- colors: 40, 40, 42, 42
		778 => x"2A2A0000",		-- colors: 42, 42, 40, 40
		779 => x"002A2A2A",		-- colors: 40, 42, 42, 42
		780 => x"2A2A2A00",		-- colors: 42, 42, 42, 40
		781 => x"002A2A2A",		-- colors: 40, 42, 42, 42
		782 => x"2A2A2A00",		-- colors: 42, 42, 42, 40
		783 => x"002A2A2A",		-- colors: 40, 42, 42, 42
		784 => x"2A2A2A00",		-- colors: 42, 42, 42, 40
		785 => x"002A2A2A",		-- colors: 40, 42, 42, 42
		786 => x"2A2A2A00",		-- colors: 42, 42, 42, 40
		787 => x"00002A2A",		-- colors: 40, 40, 42, 42
		788 => x"2A2A0000",		-- colors: 42, 42, 40, 40
		789 => x"00002A2A",		-- colors: 40, 40, 42, 42
		790 => x"2A2A0000",		-- colors: 42, 42, 40, 40
		791 => x"00000000",		-- colors: 40, 40, 40, 40
		792 => x"00000000",		-- colors: 40, 40, 40, 40
		793 => x"00000000",		-- colors: 40, 40, 40, 40
		794 => x"00000000",		-- colors: 40, 40, 40, 40
		795 => x"29292929",		-- colors: 41, 41, 41, 41
		796 => x"29292929",		-- colors: 41, 41, 41, 41
		797 => x"29292929",		-- colors: 41, 41, 41, 41
		798 => x"29292929",		-- colors: 41, 41, 41, 41
		799 => x"2B2A2A2A",		-- colors: 43, 42, 42, 42
		800 => x"2A2A2A2B",		-- colors: 42, 42, 42, 43
		801 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		802 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		803 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
		804 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
		805 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		806 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		807 => x"2B2A2A2A",		-- colors: 43, 42, 42, 42
		808 => x"2A2A2A2B",		-- colors: 42, 42, 42, 43
		809 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		810 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		811 => x"2B2A2A2A",		-- colors: 43, 42, 42, 42
		812 => x"2A2A2A2B",		-- colors: 42, 42, 42, 43
		813 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		814 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		815 => x"2B2A2A2A",		-- colors: 43, 42, 42, 42
		816 => x"2A2A2A2B",		-- colors: 42, 42, 42, 43
		817 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		818 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		819 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
		820 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
		821 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		822 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		823 => x"2B2A2A2A",		-- colors: 43, 42, 42, 42
		824 => x"2A2A2A2B",		-- colors: 42, 42, 42, 43
		825 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		826 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		827 => x"2B2A2A2A",		-- colors: 43, 42, 42, 42
		828 => x"2A2A2A2B",		-- colors: 42, 42, 42, 43
		829 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
		830 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42

				----------------------------------------------------
        6992 => x"00000016", -- pedding 
        6993 => x"00000016", -- pedding 
        6994 => x"00000016", -- pedding 
        6995 => x"00000016", -- pedding 
        6996 => x"00000016", -- pedding 
        6997 => x"00000016", -- pedding 
        6998 => x"00000016", -- pedding 
        6999 => x"00000016", -- pedding 
        7000 => x"00000016", -- pedding 
        7001 => x"00000016", -- pedding 
        7002 => x"00000016", -- pedding 
        7003 => x"00000016", -- pedding 
        7004 => x"00000016", -- pedding 
        7005 => x"00000016", -- pedding 
        7006 => x"00000016", -- pedding 
        7007 => x"00000016", -- pedding 
        7008 => x"00000016", -- pedding 
        7009 => x"00000016", -- pedding 
        7010 => x"00000016", -- pedding 
        7011 => x"00000016", -- pedding 
        7012 => x"00000016", -- pedding 
        7013 => x"00000016", -- pedding 
        7014 => x"00000016", -- pedding 
        7015 => x"00000016", -- pedding 
        7016 => x"00000016", -- pedding 
        7017 => x"00000016", -- pedding 
        7018 => x"00000016", -- pedding 
        7019 => x"00000016", -- pedding 
        7020 => x"00000016", -- pedding 
        7021 => x"00000016", -- pedding 
        7022 => x"00000016", -- pedding 
        7023 => x"00000016", -- pedding 
        7024 => x"00000016", -- pedding 
        7025 => x"00000016", -- pedding 
        7026 => x"00000016", -- pedding 
        7027 => x"00000016", -- pedding 
        7028 => x"00000016", -- pedding 
        7029 => x"00000016", -- pedding 
        7030 => x"00000016", -- pedding 
        7031 => x"00000016", -- pedding 
        7032 => x"00000016", -- pedding 
        7033 => x"00000016", -- pedding 
        7034 => x"00000016", -- pedding 
        7035 => x"00000016", -- pedding 
        7036 => x"00000016", -- pedding 
        7037 => x"00000016", -- pedding 
        7038 => x"00000016", -- pedding 
        7039 => x"00000016", -- pedding 
        7040 => x"00000016", -- pedding 
        7041 => x"00000016", -- pedding 
        7042 => x"00000016", -- pedding 
        7043 => x"00000016", -- pedding 
        7044 => x"00000016", -- pedding 
        7045 => x"00000016", -- pedding 
        7046 => x"00000016", -- pedding 
        7047 => x"00000016", -- pedding 
        7048 => x"00000016", -- pedding 
        7049 => x"00000016", -- pedding 
        7050 => x"00000016", -- pedding 
        7051 => x"00000016", -- pedding 
        7052 => x"00000016", -- pedding 
        7053 => x"00000016", -- pedding 
        7054 => x"00000016", -- pedding 
        7055 => x"00000016", -- pedding 
        7056 => x"00000016", -- pedding 
        7057 => x"00000016", -- pedding 
        7058 => x"00000016", -- pedding 
        7059 => x"00000016", -- pedding 
        7060 => x"00000016", -- pedding 
        7061 => x"00000016", -- pedding 
        7062 => x"00000016", -- pedding 
        7063 => x"00000016", -- pedding 
        7064 => x"00000016", -- pedding 
        7065 => x"00000016", -- pedding 
        7066 => x"00000016", -- pedding 
        7067 => x"00000016", -- pedding 
        7068 => x"00000016", -- pedding 
        7069 => x"00000016", -- pedding 
        7070 => x"00000016", -- pedding 
        7071 => x"00000016", -- pedding 
        7072 => x"00000016", -- pedding 
        7073 => x"00000016", -- pedding 
        7074 => x"00000016", -- pedding 
        7075 => x"00000016", -- pedding 
        7076 => x"00000016", -- pedding 
        7077 => x"00000016", -- pedding 
        7078 => x"00000016", -- pedding 
        7079 => x"00000016", -- pedding 
        7080 => x"00000016", -- pedding 
        7081 => x"00000016", -- pedding 
        7082 => x"00000016", -- pedding 
        7083 => x"00000016", -- pedding 
        7084 => x"00000016", -- pedding 
        7085 => x"00000016", -- pedding 
        7086 => x"00000016", -- pedding 
        7087 => x"00000016", -- pedding 
        7088 => x"00000016", -- pedding 
        7089 => x"00000016", -- pedding 
        7090 => x"00000016", -- pedding 
        7091 => x"00000016", -- pedding 
        7092 => x"00000016", -- pedding 
        7093 => x"00000016", -- pedding 
        7094 => x"00000016", -- pedding 
        7095 => x"00000016", -- pedding 
        7096 => x"00000016", -- pedding 
        7097 => x"00000016", -- pedding 
        7098 => x"00000016", -- pedding 
        7099 => x"00000016", -- pedding 
        7100 => x"00000016", -- pedding 
        7101 => x"00000016", -- pedding 
        7102 => x"00000016", -- pedding 
        7103 => x"00000016", -- pedding 
        7104 => x"00000016", -- pedding 
        7105 => x"00000016", -- pedding 
        7106 => x"00000016", -- pedding 
        7107 => x"00000016", -- pedding 
        7108 => x"00000016", -- pedding 
        7109 => x"00000016", -- pedding 
        7110 => x"00000016", -- pedding 
        7111 => x"00000016", -- pedding 
        7112 => x"00000016", -- pedding 
        7113 => x"00000016", -- pedding 
        7114 => x"00000016", -- pedding 
        7115 => x"00000016", -- pedding 
        7116 => x"00000016", -- pedding 
        7117 => x"00000016", -- pedding 
        7118 => x"00000016", -- pedding 
        7119 => x"00000016", -- pedding 
        7120 => x"00000016", -- pedding 
        7121 => x"00000016", -- pedding 
        7122 => x"00000016", -- pedding 
        7123 => x"00000016", -- pedding 
        7124 => x"00000016", -- header 
        7125 => x"00000016", -- header 
        7126 => x"00000016", -- header 
        7127 => x"00000016", -- header 
        7128 => x"00000016", -- header 
        7129 => x"00000016", -- header 
        7130 => x"00000016", -- header 
        7131 => x"00000016", -- header 
        7132 => x"00000016", -- header 
        7133 => x"00000016", -- header 
        7134 => x"00000016", -- header 
        7135 => x"00000016", -- header 
        7136 => x"00000016", -- header 
        7137 => x"00000016", -- header 
        7138 => x"00000016", -- header 
        7139 => x"00000016", -- header 
        7140 => x"00000016", -- pedding 
        7141 => x"00000016", -- pedding 
        7142 => x"00000016", -- pedding 
        7143 => x"00000016", -- pedding 
        7144 => x"00000016", -- pedding 
        7145 => x"00000016", -- pedding 
        7146 => x"00000016", -- pedding 
        7147 => x"00000016", -- pedding 
        7148 => x"00000016", -- pedding 
        7149 => x"00000016", -- pedding 
        7150 => x"00000016", -- pedding 
        7151 => x"00000016", -- pedding 
        7152 => x"00000016", -- pedding 
        7153 => x"00000016", -- pedding 
        7154 => x"00000016", -- pedding 
        7155 => x"00000016", -- pedding 
        7156 => x"00000016", -- pedding 
        7157 => x"00000016", -- pedding 
        7158 => x"00000016", -- pedding 
        7159 => x"00000016", -- pedding 
        7160 => x"00000016", -- pedding 
        7161 => x"00000016", -- pedding 
        7162 => x"00000016", -- pedding 
        7163 => x"00000016", -- pedding 
        7164 => x"00000016", -- header 
        7165 => x"00000016", -- header 
        7166 => x"00000016", -- header 
        7167 => x"00000016", -- header 
        7168 => x"00000016", -- header 
        7169 => x"00000016", -- header 
        7170 => x"00000016", -- header 
        7171 => x"00000016", -- header 
        7172 => x"00000016", -- header 
        7173 => x"00000016", -- header 
        7174 => x"00000016", -- header 
        7175 => x"00000016", -- header 
        7176 => x"00000016", -- header 
        7177 => x"00000016", -- header 
        7178 => x"00000016", -- header 
        7179 => x"00000016", -- header 
        7180 => x"00000016", -- pedding 
        7181 => x"00000016", -- pedding 
        7182 => x"00000016", -- pedding 
        7183 => x"00000016", -- pedding 
        7184 => x"00000016", -- pedding 
        7185 => x"00000016", -- pedding 
        7186 => x"00000016", -- pedding 
        7187 => x"00000016", -- pedding 
        7188 => x"00000016", -- pedding 
        7189 => x"00000016", -- pedding 
        7190 => x"00000016", -- pedding 
        7191 => x"00000016", -- pedding 
        7192 => x"00000016", -- pedding 
        7193 => x"00000016", -- pedding 
        7194 => x"00000016", -- pedding 
        7195 => x"00000016", -- pedding 
        7196 => x"00000016", -- pedding 
        7197 => x"00000016", -- pedding 
        7198 => x"00000016", -- pedding 
        7199 => x"00000016", -- pedding 
        7200 => x"00000016", -- pedding 
        7201 => x"00000016", -- pedding 
        7202 => x"00000016", -- pedding 
        7203 => x"00000016", -- pedding 
        7204 => x"00000016", -- header 
        7205 => x"00000016", -- header 
        7206 => x"00000016", -- header 
        7207 => x"00000016", -- header 
        7208 => x"00000016", -- header 
        7209 => x"00000016", -- header 
        7210 => x"00000016", -- header 
        7211 => x"00000016", -- header 
        7212 => x"00000016", -- header 
        7213 => x"00000016", -- header 
        7214 => x"00000016", -- header 
        7215 => x"00000016", -- header 
        7216 => x"00000016", -- header 
        7217 => x"00000016", -- header 
        7218 => x"00000016", -- header 
        7219 => x"00000016", -- header 
        7220 => x"00000016", -- pedding 
        7221 => x"00000016", -- pedding 
        7222 => x"00000016", -- pedding 
        7223 => x"00000016", -- pedding 
        7224 => x"00000016", -- pedding 
        7225 => x"00000016", -- pedding 
        7226 => x"00000016", -- pedding 
        7227 => x"00000016", -- pedding 
        7228 => x"00000016", -- pedding 
        7229 => x"00000016", -- pedding 
        7230 => x"00000016", -- pedding 
        7231 => x"00000016", -- pedding 
        7232 => x"00000016", -- pedding 
        7233 => x"00000016", -- pedding 
        7234 => x"00000016", -- pedding 
        7235 => x"00000016", -- pedding 
        7236 => x"00000016", -- pedding 
        7237 => x"00000016", -- pedding 
        7238 => x"00000016", -- pedding 
        7239 => x"00000016", -- pedding 
        7240 => x"00000016", -- pedding 
        7241 => x"00000016", -- pedding 
        7242 => x"00000016", -- pedding 
        7243 => x"00000016", -- pedding 
        7244 => x"00000016", -- header 
        7245 => x"00000016", -- header 
        7246 => x"00000016", -- header 
        7247 => x"00000016", -- header 
        7248 => x"00000016", -- header 
        7249 => x"00000016", -- header 
        7250 => x"00000016", -- header 
        7251 => x"00000016", -- header 
        7252 => x"00000016", -- header 
        7253 => x"00000016", -- header 
        7254 => x"00000016", -- header 
        7255 => x"00000016", -- header 
        7256 => x"00000016", -- header 
        7257 => x"00000016", -- header 
        7258 => x"00000016", -- header 
        7259 => x"00000016", -- header 
        7260 => x"00000016", -- pedding 
        7261 => x"00000016", -- pedding 
        7262 => x"00000016", -- pedding 
        7263 => x"00000016", -- pedding 
        7264 => x"00000016", -- pedding 
        7265 => x"00000016", -- pedding 
        7266 => x"00000016", -- pedding 
        7267 => x"00000016", -- pedding 
        7268 => x"00000016", -- pedding 
        7269 => x"00000016", -- pedding 
        7270 => x"00000016", -- pedding 
        7271 => x"00000016", -- pedding 
        7272 => x"00000016", -- pedding 
        7273 => x"00000016", -- pedding 
        7274 => x"00000016", -- pedding 
        7275 => x"00000016", -- pedding 
        7276 => x"00000016", -- pedding 
        7277 => x"00000016", -- pedding 
        7278 => x"00000016", -- pedding 
        7279 => x"00000016", -- pedding 
        7280 => x"00000016", -- pedding 
        7281 => x"00000016", -- pedding 
        7282 => x"00000016", -- pedding 
        7283 => x"00000016", -- pedding 
        7284 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7285 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7286 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7287 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7288 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7289 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7290 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7291 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7292 => x"00000001", -- z: 0 rot: 0 ptr: 319
        7293 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7294 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7295 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7296 => x"00000001", -- z: 0 rot: 0 ptr: 319
        7297 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7298 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7299 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7300 => x"00000016", -- pedding 
        7301 => x"00000016", -- pedding 
        7302 => x"00000016", -- pedding 
        7303 => x"00000016", -- pedding 
        7304 => x"00000016", -- pedding 
        7305 => x"00000016", -- pedding 
        7306 => x"00000016", -- pedding 
        7307 => x"00000016", -- pedding 
        7308 => x"00000016", -- pedding 
        7309 => x"00000016", -- pedding 
        7310 => x"00000016", -- pedding 
        7311 => x"00000016", -- pedding 
        7312 => x"00000016", -- pedding 
        7313 => x"00000016", -- pedding 
        7314 => x"00000016", -- pedding 
        7315 => x"00000016", -- pedding 
        7316 => x"00000016", -- pedding 
        7317 => x"00000016", -- pedding 
        7318 => x"00000016", -- pedding 
        7319 => x"00000016", -- pedding 
        7320 => x"00000016", -- pedding 
        7321 => x"00000016", -- pedding 
        7322 => x"00000016", -- pedding 
        7323 => x"00000016", -- pedding 
        7324 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7325 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7326 => x"00000003", -- z: 0 rot: 0 ptr: 447
        7327 => x"00000005", -- z: 0 rot: 0 ptr: 575
        7328 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7329 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7330 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7331 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7332 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7333 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7334 => x"00000001", -- z: 0 rot: 0 ptr: 319
        7335 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7336 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7337 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7338 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7339 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7340 => x"00000016", -- pedding 
        7341 => x"00000016", -- pedding 
        7342 => x"00000016", -- pedding 
        7343 => x"00000016", -- pedding 
        7344 => x"00000016", -- pedding 
        7345 => x"00000016", -- pedding 
        7346 => x"00000016", -- pedding 
        7347 => x"00000016", -- pedding 
        7348 => x"00000016", -- pedding 
        7349 => x"00000016", -- pedding 
        7350 => x"00000016", -- pedding 
        7351 => x"00000016", -- pedding 
        7352 => x"00000016", -- pedding 
        7353 => x"00000016", -- pedding 
        7354 => x"00000016", -- pedding 
        7355 => x"00000016", -- pedding 
        7356 => x"00000016", -- pedding 
        7357 => x"00000016", -- pedding 
        7358 => x"00000016", -- pedding 
        7359 => x"00000016", -- pedding 
        7360 => x"00000016", -- pedding 
        7361 => x"00000016", -- pedding 
        7362 => x"00000016", -- pedding 
        7363 => x"00000016", -- pedding 
        7364 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7365 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7366 => x"00000015", -- z: 0 rot: 0 ptr: 831
        7367 => x"00000017", -- z: 0 rot: 0 ptr: 959
        7368 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7369 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7370 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7371 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7372 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7373 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7374 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7375 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7376 => x"00000001", -- z: 0 rot: 0 ptr: 319
        7377 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7378 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7379 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7380 => x"00000016", -- pedding 
        7381 => x"00000016", -- pedding 
        7382 => x"00000016", -- pedding 
        7383 => x"00000016", -- pedding 
        7384 => x"00000016", -- pedding 
        7385 => x"00000016", -- pedding 
        7386 => x"00000016", -- pedding 
        7387 => x"00000016", -- pedding 
        7388 => x"00000016", -- pedding 
        7389 => x"00000016", -- pedding 
        7390 => x"00000016", -- pedding 
        7391 => x"00000016", -- pedding 
        7392 => x"00000016", -- pedding 
        7393 => x"00000016", -- pedding 
        7394 => x"00000016", -- pedding 
        7395 => x"00000016", -- pedding 
        7396 => x"00000016", -- pedding 
        7397 => x"00000016", -- pedding 
        7398 => x"00000016", -- pedding 
        7399 => x"00000016", -- pedding 
        7400 => x"00000016", -- pedding 
        7401 => x"00000016", -- pedding 
        7402 => x"00000016", -- pedding 
        7403 => x"00000016", -- pedding 
        7404 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7405 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7406 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7407 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7408 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7409 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7410 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7411 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7412 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7413 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7414 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7415 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7416 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7417 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7418 => x"00000024", -- z: 0 rot: 0 ptr: 1023
        7419 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7420 => x"00000016", -- pedding 
        7421 => x"00000016", -- pedding 
        7422 => x"00000016", -- pedding 
        7423 => x"00000016", -- pedding 
        7424 => x"00000016", -- pedding 
        7425 => x"00000016", -- pedding 
        7426 => x"00000016", -- pedding 
        7427 => x"00000016", -- pedding 
        7428 => x"00000016", -- pedding 
        7429 => x"00000016", -- pedding 
        7430 => x"00000016", -- pedding 
        7431 => x"00000016", -- pedding 
        7432 => x"00000016", -- pedding 
        7433 => x"00000016", -- pedding 
        7434 => x"00000016", -- pedding 
        7435 => x"00000016", -- pedding 
        7436 => x"00000016", -- pedding 
        7437 => x"00000016", -- pedding 
        7438 => x"00000016", -- pedding 
        7439 => x"00000016", -- pedding 
        7440 => x"00000016", -- pedding 
        7441 => x"00000016", -- pedding 
        7442 => x"00000016", -- pedding 
        7443 => x"00000016", -- pedding 
        7444 => x"00000025", -- z: 0 rot: 0 ptr: 1087
        7445 => x"00000025", -- z: 0 rot: 0 ptr: 1087
        7446 => x"00000025", -- z: 0 rot: 0 ptr: 1087
        7447 => x"00000025", -- z: 0 rot: 0 ptr: 1087
        7448 => x"00000025", -- z: 0 rot: 0 ptr: 1087
        7449 => x"00000025", -- z: 0 rot: 0 ptr: 1087
        7450 => x"00000025", -- z: 0 rot: 0 ptr: 1087
        7451 => x"00000025", -- z: 0 rot: 0 ptr: 1087
        7452 => x"00000025", -- z: 0 rot: 0 ptr: 1087
        7453 => x"00000025", -- z: 0 rot: 0 ptr: 1087
        7454 => x"00000025", -- z: 0 rot: 0 ptr: 1087
        7455 => x"00000025", -- z: 0 rot: 0 ptr: 1087
        7456 => x"00000025", -- z: 0 rot: 0 ptr: 1087
        7457 => x"00000025", -- z: 0 rot: 0 ptr: 1087
        7458 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7459 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7460 => x"00000016", -- pedding 
        7461 => x"00000016", -- pedding 
        7462 => x"00000016", -- pedding 
        7463 => x"00000016", -- pedding 
        7464 => x"00000016", -- pedding 
        7465 => x"00000016", -- pedding 
        7466 => x"00000016", -- pedding 
        7467 => x"00000016", -- pedding 
        7468 => x"00000016", -- pedding 
        7469 => x"00000016", -- pedding 
        7470 => x"00000016", -- pedding 
        7471 => x"00000016", -- pedding 
        7472 => x"00000016", -- pedding 
        7473 => x"00000016", -- pedding 
        7474 => x"00000016", -- pedding 
        7475 => x"00000016", -- pedding 
        7476 => x"00000016", -- pedding 
        7477 => x"00000016", -- pedding 
        7478 => x"00000016", -- pedding 
        7479 => x"00000016", -- pedding 
        7480 => x"00000016", -- pedding 
        7481 => x"00000016", -- pedding 
        7482 => x"00000016", -- pedding 
        7483 => x"00000016", -- pedding 
        7484 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7485 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7486 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7487 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7488 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7489 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7490 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7491 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7492 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7493 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7494 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7495 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7496 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7497 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7498 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7499 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7500 => x"00000016", -- pedding 
        7501 => x"00000016", -- pedding 
        7502 => x"00000016", -- pedding 
        7503 => x"00000016", -- pedding 
        7504 => x"00000016", -- pedding 
        7505 => x"00000016", -- pedding 
        7506 => x"00000016", -- pedding 
        7507 => x"00000016", -- pedding 
        7508 => x"00000016", -- pedding 
        7509 => x"00000016", -- pedding 
        7510 => x"00000016", -- pedding 
        7511 => x"00000016", -- pedding 
        7512 => x"00000016", -- pedding 
        7513 => x"00000016", -- pedding 
        7514 => x"00000016", -- pedding 
        7515 => x"00000016", -- pedding 
        7516 => x"00000016", -- pedding 
        7517 => x"00000016", -- pedding 
        7518 => x"00000016", -- pedding 
        7519 => x"00000016", -- pedding 
        7520 => x"00000016", -- pedding 
        7521 => x"00000016", -- pedding 
        7522 => x"00000016", -- pedding 
        7523 => x"00000016", -- pedding 
        7524 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7525 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7526 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7527 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7528 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7529 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7530 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7531 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7532 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7533 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7534 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7535 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7536 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7537 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7538 => x"00000013", -- z: 0 rot: 0 ptr: 703
        7539 => x"00000013", -- z: 0 rot: 0 ptr: 703
        7540 => x"00000016", -- pedding 
        7541 => x"00000016", -- pedding 
        7542 => x"00000016", -- pedding 
        7543 => x"00000016", -- pedding 
        7544 => x"00000016", -- pedding 
        7545 => x"00000016", -- pedding 
        7546 => x"00000016", -- pedding 
        7547 => x"00000016", -- pedding 
        7548 => x"00000016", -- pedding 
        7549 => x"00000016", -- pedding 
        7550 => x"00000016", -- pedding 
        7551 => x"00000016", -- pedding 
        7552 => x"00000016", -- pedding 
        7553 => x"00000016", -- pedding 
        7554 => x"00000016", -- pedding 
        7555 => x"00000016", -- pedding 
        7556 => x"00000016", -- pedding 
        7557 => x"00000016", -- pedding 
        7558 => x"00000016", -- pedding 
        7559 => x"00000016", -- pedding 
        7560 => x"00000016", -- pedding 
        7561 => x"00000016", -- pedding 
        7562 => x"00000016", -- pedding 
        7563 => x"00000016", -- pedding 
        7564 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7565 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7566 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7567 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7568 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7569 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7570 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7571 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7572 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7573 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7574 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7575 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7576 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7577 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7578 => x"00000013", -- z: 0 rot: 0 ptr: 703
        7579 => x"00000013", -- z: 0 rot: 0 ptr: 703
        7580 => x"00000016", -- pedding 
        7581 => x"00000016", -- pedding 
        7582 => x"00000016", -- pedding 
        7583 => x"00000016", -- pedding 
        7584 => x"00000016", -- pedding 
        7585 => x"00000016", -- pedding 
        7586 => x"00000016", -- pedding 
        7587 => x"00000016", -- pedding 
        7588 => x"00000016", -- pedding 
        7589 => x"00000016", -- pedding 
        7590 => x"00000016", -- pedding 
        7591 => x"00000016", -- pedding 
        7592 => x"00000016", -- pedding 
        7593 => x"00000016", -- pedding 
        7594 => x"00000016", -- pedding 
        7595 => x"00000016", -- pedding 
        7596 => x"00000016", -- pedding 
        7597 => x"00000016", -- pedding 
        7598 => x"00000016", -- pedding 
        7599 => x"00000016", -- pedding 
        7600 => x"00000016", -- pedding 
        7601 => x"00000016", -- pedding 
        7602 => x"00000016", -- pedding 
        7603 => x"00000016", -- pedding 
        7604 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7605 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7606 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7607 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7608 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7609 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7610 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7611 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7612 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7613 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7614 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7615 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7616 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7617 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7618 => x"00000013", -- z: 0 rot: 0 ptr: 703
        7619 => x"00000013", -- z: 0 rot: 0 ptr: 703
        7620 => x"00000016", -- pedding 
        7621 => x"00000016", -- pedding 
        7622 => x"00000016", -- pedding 
        7623 => x"00000016", -- pedding 
        7624 => x"00000016", -- pedding 
        7625 => x"00000016", -- pedding 
        7626 => x"00000016", -- pedding 
        7627 => x"00000016", -- pedding 
        7628 => x"00000016", -- pedding 
        7629 => x"00000016", -- pedding 
        7630 => x"00000016", -- pedding 
        7631 => x"00000016", -- pedding 
        7632 => x"00000016", -- pedding 
        7633 => x"00000016", -- pedding 
        7634 => x"00000016", -- pedding 
        7635 => x"00000016", -- pedding 
        7636 => x"00000016", -- pedding 
        7637 => x"00000016", -- pedding 
        7638 => x"00000016", -- pedding 
        7639 => x"00000016", -- pedding 
        7640 => x"00000016", -- pedding 
        7641 => x"00000016", -- pedding 
        7642 => x"00000016", -- pedding 
        7643 => x"00000016", -- pedding 
        7644 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7645 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7646 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7647 => x"00000092", -- z: 0 rot: 0 ptr: 3455
        7648 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7649 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7650 => x"00000092", -- z: 0 rot: 0 ptr: 3455
        7651 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7652 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7653 => x"00000092", -- z: 0 rot: 0 ptr: 3455
        7654 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7655 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7656 => x"00000092", -- z: 0 rot: 0 ptr: 3455
        7657 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7658 => x"00000013", -- z: 0 rot: 0 ptr: 703
        7659 => x"00000013", -- z: 0 rot: 0 ptr: 703
        7660 => x"00000016", -- pedding 
        7661 => x"00000016", -- pedding 
        7662 => x"00000016", -- pedding 
        7663 => x"00000016", -- pedding 
        7664 => x"00000016", -- pedding 
        7665 => x"00000016", -- pedding 
        7666 => x"00000016", -- pedding 
        7667 => x"00000016", -- pedding 
        7668 => x"00000016", -- pedding 
        7669 => x"00000016", -- pedding 
        7670 => x"00000016", -- pedding 
        7671 => x"00000016", -- pedding 
        7672 => x"00000016", -- pedding 
        7673 => x"00000016", -- pedding 
        7674 => x"00000016", -- pedding 
        7675 => x"00000016", -- pedding 
        7676 => x"00000016", -- pedding 
        7677 => x"00000016", -- pedding 
        7678 => x"00000016", -- pedding 
        7679 => x"00000016", -- pedding 
        7680 => x"00000016", -- pedding 
        7681 => x"00000016", -- pedding 
        7682 => x"00000016", -- pedding 
        7683 => x"00000016", -- pedding 
        7684 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7685 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7686 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7687 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7688 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7689 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7690 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7691 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7692 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7693 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7694 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7695 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7696 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7697 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7698 => x"00000013", -- z: 0 rot: 0 ptr: 703
        7699 => x"00000013", -- z: 0 rot: 0 ptr: 703
        7700 => x"00000016", -- pedding 
        7701 => x"00000016", -- pedding 
        7702 => x"00000016", -- pedding 
        7703 => x"00000016", -- pedding 
        7704 => x"00000016", -- pedding 
        7705 => x"00000016", -- pedding 
        7706 => x"00000016", -- pedding 
        7707 => x"00000016", -- pedding 
        7708 => x"00000016", -- pedding 
        7709 => x"00000016", -- pedding 
        7710 => x"00000016", -- pedding 
        7711 => x"00000016", -- pedding 
        7712 => x"00000016", -- pedding 
        7713 => x"00000016", -- pedding 
        7714 => x"00000016", -- pedding 
        7715 => x"00000016", -- pedding 
        7716 => x"00000016", -- pedding 
        7717 => x"00000016", -- pedding 
        7718 => x"00000016", -- pedding 
        7719 => x"00000016", -- pedding 
        7720 => x"00000016", -- pedding 
        7721 => x"00000016", -- pedding 
        7722 => x"00000016", -- pedding 
        7723 => x"00000016", -- pedding 
        7724 => x"00000016", -- pedding 
        7725 => x"00000016", -- pedding 
        7726 => x"00000016", -- pedding 
        7727 => x"00000016", -- pedding 
        7728 => x"00000016", -- pedding 
        7729 => x"00000016", -- pedding 
        7730 => x"00000016", -- pedding 
        7731 => x"00000016", -- pedding 
        7732 => x"00000016", -- pedding 
        7733 => x"00000016", -- pedding 
        7734 => x"00000016", -- pedding 
        7735 => x"00000016", -- pedding 
        7736 => x"00000016", -- pedding 
        7737 => x"00000016", -- pedding 
        7738 => x"00000016", -- pedding 
        7739 => x"00000016", -- pedding 
        7740 => x"00000016", -- pedding 
        7741 => x"00000016", -- pedding 
        7742 => x"00000016", -- pedding 
        7743 => x"00000016", -- pedding 
        7744 => x"00000016", -- pedding 
        7745 => x"00000016", -- pedding 
        7746 => x"00000016", -- pedding 
        7747 => x"00000016", -- pedding 
        7748 => x"00000016", -- pedding 
        7749 => x"00000016", -- pedding 
        7750 => x"00000016", -- pedding 
        7751 => x"00000016", -- pedding 
        7752 => x"00000016", -- pedding 
        7753 => x"00000016", -- pedding 
        7754 => x"00000016", -- pedding 
        7755 => x"00000016", -- pedding 
        7756 => x"00000016", -- pedding 
        7757 => x"00000016", -- pedding 
        7758 => x"00000016", -- pedding 
        7759 => x"00000016", -- pedding 
        7760 => x"00000016", -- pedding 
        7761 => x"00000016", -- pedding 
        7762 => x"00000016", -- pedding 
        7763 => x"00000016", -- pedding 
        7764 => x"00000016", -- pedding 
        7765 => x"00000016", -- pedding 
        7766 => x"00000016", -- pedding 
        7767 => x"00000016", -- pedding 
        7768 => x"00000016", -- pedding 
        7769 => x"00000016", -- pedding 
        7770 => x"00000016", -- pedding 
        7771 => x"00000016", -- pedding 
        7772 => x"00000016", -- pedding 
        7773 => x"00000016", -- pedding 
        7774 => x"00000016", -- pedding 
        7775 => x"00000016", -- pedding 
        7776 => x"00000016", -- pedding 
        7777 => x"00000016", -- pedding 
        7778 => x"00000016", -- pedding 
        7779 => x"00000016", -- pedding 
        7780 => x"00000016", -- pedding 
        7781 => x"00000016", -- pedding 
        7782 => x"00000016", -- pedding 
        7783 => x"00000016", -- pedding 
        7784 => x"00000016", -- pedding 
        7785 => x"00000016", -- pedding 
        7786 => x"00000016", -- pedding 
        7787 => x"00000016", -- pedding 
        7788 => x"00000016", -- pedding 
        7789 => x"00000016", -- pedding 
        7790 => x"00000016", -- pedding 
        7791 => x"00000016", -- pedding 
        7792 => x"00000016", -- pedding 
        7793 => x"00000016", -- pedding 
        7794 => x"00000016", -- pedding 
        7795 => x"00000016", -- pedding 
        7796 => x"00000016", -- pedding 
        7797 => x"00000016", -- pedding 
        7798 => x"00000016", -- pedding 
        7799 => x"00000016", -- pedding 
        7800 => x"00000016", -- pedding 
        7801 => x"00000016", -- pedding 
        7802 => x"00000016", -- pedding 
        7803 => x"00000016", -- pedding 
        7804 => x"00000016", -- pedding 
        7805 => x"00000016", -- pedding 
        7806 => x"00000016", -- pedding 
        7807 => x"00000016", -- pedding 
        7808 => x"00000016", -- pedding 
        7809 => x"00000016", -- pedding 
        7810 => x"00000016", -- pedding 
        7811 => x"00000016", -- pedding 
        7812 => x"00000016", -- pedding 
        7813 => x"00000016", -- pedding 
        7814 => x"00000016", -- pedding 
        7815 => x"00000016", -- pedding 
        7816 => x"00000016", -- pedding 
        7817 => x"00000016", -- pedding 
        7818 => x"00000016", -- pedding 
        7819 => x"00000016", -- pedding 
        7820 => x"00000016", -- pedding 
        7821 => x"00000016", -- pedding 
        7822 => x"00000016", -- pedding 
        7823 => x"00000016", -- pedding 
        7824 => x"00000016", -- pedding 
        7825 => x"00000016", -- pedding 
        7826 => x"00000016", -- pedding 
        7827 => x"00000016", -- pedding 
        7828 => x"00000016", -- pedding 
        7829 => x"00000016", -- pedding 
        7830 => x"00000016", -- pedding 
        7831 => x"00000016", -- pedding 
        7832 => x"00000016", -- pedding 
        7833 => x"00000016", -- pedding 
        7834 => x"00000016", -- pedding 
        7835 => x"00000016", -- pedding 
        7836 => x"00000016", -- pedding 
        7837 => x"00000016", -- pedding 
        7838 => x"00000016", -- pedding 
        7839 => x"00000016", -- pedding 
        7840 => x"00000016", -- pedding 
        7841 => x"00000016", -- pedding 
        7842 => x"00000016", -- pedding 
        7843 => x"00000016", -- pedding 
        7844 => x"00000016", -- pedding 
        7845 => x"00000016", -- pedding 
        7846 => x"00000016", -- pedding 
        7847 => x"00000016", -- pedding 
        7848 => x"00000016", -- pedding 
        7849 => x"00000016", -- pedding 
        7850 => x"00000016", -- pedding 
        7851 => x"00000016", -- pedding 
        7852 => x"00000016", -- pedding 
        7853 => x"00000016", -- pedding 
        7854 => x"00000016", -- pedding 
        7855 => x"00000016", -- pedding 
        7856 => x"00000016", -- pedding 
        7857 => x"00000016", -- pedding 
        7858 => x"00000016", -- pedding 
        7859 => x"00000016", -- pedding 
        7860 => x"00000016", -- pedding 
        7861 => x"00000016", -- pedding 
        7862 => x"00000016", -- pedding 
        7863 => x"00000016", -- pedding 
        7864 => x"00000016", -- pedding 
        7865 => x"00000016", -- pedding 
        7866 => x"00000016", -- pedding 
        7867 => x"00000016", -- pedding 
        7868 => x"00000016", -- pedding 
        7869 => x"00000016", -- pedding 
        7870 => x"00000016", -- pedding 
        7871 => x"00000016", -- pedding 
        7872 => x"00000016", -- pedding 
        7873 => x"00000016", -- pedding 
        7874 => x"00000016", -- pedding 
        7875 => x"00000016", -- pedding 
        7876 => x"00000016", -- pedding 
        7877 => x"00000016", -- pedding 
        7878 => x"00000016", -- pedding 
        7879 => x"00000016", -- pedding 
        7880 => x"00000016", -- pedding 
        7881 => x"00000016", -- pedding 
        7882 => x"00000016", -- pedding 
        7883 => x"00000016", -- pedding 
        7884 => x"00000016", -- pedding 
        7885 => x"00000016", -- pedding 
        7886 => x"00000016", -- pedding 
        7887 => x"00000016", -- pedding 
        7888 => x"00000016", -- pedding 
        7889 => x"00000016", -- pedding 
        7890 => x"00000016", -- pedding 
        7891 => x"00000016", -- pedding 
        7892 => x"00000016", -- pedding 
        7893 => x"00000016", -- pedding 
        7894 => x"00000016", -- pedding 
        7895 => x"00000016", -- pedding 
        7896 => x"00000016", -- pedding 
        7897 => x"00000016", -- pedding 
        7898 => x"00000016", -- pedding 
        7899 => x"00000016", -- pedding 
        7900 => x"00000016", -- pedding 
        7901 => x"00000016", -- pedding 
        7902 => x"00000016", -- pedding 
        7903 => x"00000016", -- pedding 
        7904 => x"00000016", -- pedding 
        7905 => x"00000016", -- pedding 
        7906 => x"00000016", -- pedding 
        7907 => x"00000016", -- pedding 
        7908 => x"00000016", -- pedding 
        7909 => x"00000016", -- pedding 
        7910 => x"00000016", -- pedding 
        7911 => x"00000016", -- pedding 
        7912 => x"00000016", -- pedding 
        7913 => x"00000016", -- pedding 
        7914 => x"00000016", -- pedding 
        7915 => x"00000016", -- pedding 
        7916 => x"00000016", -- pedding 
        7917 => x"00000016", -- pedding 
        7918 => x"00000016", -- pedding 
        7919 => x"00000016", -- pedding 
        7920 => x"00000016", -- pedding 
        7921 => x"00000016", -- pedding 
        7922 => x"00000016", -- pedding 
        7923 => x"00000016", -- pedding 
        7924 => x"00000016", -- pedding 
        7925 => x"00000016", -- pedding 
        7926 => x"00000016", -- pedding 
        7927 => x"00000016", -- pedding 
        7928 => x"00000016", -- pedding 
        7929 => x"00000016", -- pedding 
        7930 => x"00000016", -- pedding 
        7931 => x"00000016", -- pedding 
        7932 => x"00000016", -- pedding 
        7933 => x"00000016", -- pedding 
        7934 => x"00000016", -- pedding 
        7935 => x"00000016", -- pedding 
        7936 => x"00000016", -- pedding 
        7937 => x"00000016", -- pedding 
        7938 => x"00000016", -- pedding 
        7939 => x"00000016", -- pedding 
        7940 => x"00000016", -- pedding 
        7941 => x"00000016", -- pedding 
        7942 => x"00000016", -- pedding 
        7943 => x"00000016", -- pedding 
        7944 => x"00000016", -- pedding 
        7945 => x"00000016", -- pedding 
        7946 => x"00000016", -- pedding 
        7947 => x"00000016", -- pedding 
        7948 => x"00000016", -- pedding 
        7949 => x"00000016", -- pedding 
        7950 => x"00000016", -- pedding 
        7951 => x"00000016", -- pedding 
        7952 => x"00000016", -- pedding 
        7953 => x"00000016", -- pedding 
        7954 => x"00000016", -- pedding 
        7955 => x"00000016", -- pedding 
        7956 => x"00000016", -- pedding 
        7957 => x"00000016", -- pedding 
        7958 => x"00000016", -- pedding 
        7959 => x"00000016", -- pedding 
        7960 => x"00000016", -- pedding 
        7961 => x"00000016", -- pedding 
        7962 => x"00000016", -- pedding 
        7963 => x"00000016", -- pedding 
        7964 => x"00000016", -- pedding 
        7965 => x"00000016", -- pedding 
        7966 => x"00000016", -- pedding 
        7967 => x"00000016", -- pedding 
        7968 => x"00000016", -- pedding 
        7969 => x"00000016", -- pedding 
        7970 => x"00000016", -- pedding 
        7971 => x"00000016", -- pedding 
        7972 => x"00000016", -- pedding 
        7973 => x"00000016", -- pedding 
        7974 => x"00000016", -- pedding 
        7975 => x"00000016", -- pedding 
        7976 => x"00000016", -- pedding 
        7977 => x"00000016", -- pedding 
        7978 => x"00000016", -- pedding 
        7979 => x"00000016", -- pedding 
        7980 => x"00000016", -- pedding 
        7981 => x"00000016", -- pedding 
        7982 => x"00000016", -- pedding 
        7983 => x"00000016", -- pedding 
        7984 => x"00000016", -- pedding 
        7985 => x"00000016", -- pedding 
        7986 => x"00000016", -- pedding 
        7987 => x"00000016", -- pedding 
        7988 => x"00000016", -- pedding 
        7989 => x"00000016", -- pedding 
        7990 => x"00000016", -- pedding 
        7991 => x"00000016", -- pedding 
        7992 => x"00000016", -- pedding 
        7993 => x"00000016", -- pedding 
        7994 => x"00000016", -- pedding 
        7995 => x"00000016", -- pedding 
        7996 => x"00000016", -- pedding 
        7997 => x"00000016", -- pedding 
        7998 => x"00000016", -- pedding 
        7999 => x"00000016", -- pedding 
        8000 => x"00000016", -- pedding 
        8001 => x"00000016", -- pedding 
        8002 => x"00000016", -- pedding 
        8003 => x"00000016", -- pedding 
        8004 => x"00000016", -- pedding 
        8005 => x"00000016", -- pedding 
        8006 => x"00000016", -- pedding 
        8007 => x"00000016", -- pedding 
        8008 => x"00000016", -- pedding 
        8009 => x"00000016", -- pedding 
        8010 => x"00000016", -- pedding 
        8011 => x"00000016", -- pedding 
        8012 => x"00000016", -- pedding 
        8013 => x"00000016", -- pedding 
        8014 => x"00000016", -- pedding 
        8015 => x"00000016", -- pedding 
        8016 => x"00000016", -- pedding 
        8017 => x"00000016", -- pedding 
        8018 => x"00000016", -- pedding 
        8019 => x"00000016", -- pedding 
        8020 => x"00000016", -- pedding 
        8021 => x"00000016", -- pedding 
        8022 => x"00000016", -- pedding 
        8023 => x"00000016", -- pedding 
        8024 => x"00000016", -- pedding 
        8025 => x"00000016", -- pedding 
        8026 => x"00000016", -- pedding 
        8027 => x"00000016", -- pedding 
        8028 => x"00000016", -- pedding 
        8029 => x"00000016", -- pedding 
        8030 => x"00000016", -- pedding 
        8031 => x"00000016", -- pedding 
        8032 => x"00000016", -- pedding 
        8033 => x"00000016", -- pedding 
        8034 => x"00000016", -- pedding 
        8035 => x"00000016", -- pedding 
        8036 => x"00000016", -- pedding 
        8037 => x"00000016", -- pedding 
        8038 => x"00000016", -- pedding 
        8039 => x"00000016", -- pedding 
        8040 => x"00000016", -- pedding 
        8041 => x"00000016", -- pedding 
        8042 => x"00000016", -- pedding 
        8043 => x"00000016", -- pedding 
        8044 => x"00000016", -- pedding 
        8045 => x"00000016", -- pedding 
        8046 => x"00000016", -- pedding 
        8047 => x"00000016", -- pedding 
        8048 => x"00000016", -- pedding 
        8049 => x"00000016", -- pedding 
        8050 => x"00000016", -- pedding 
        8051 => x"00000016", -- pedding 
        8052 => x"00000016", -- pedding 
        8053 => x"00000016", -- pedding 
        8054 => x"00000016", -- pedding 
        8055 => x"00000016", -- pedding 
        8056 => x"00000016", -- pedding 
        8057 => x"00000016", -- pedding 
        8058 => x"00000016", -- pedding 
        8059 => x"00000016", -- pedding 
        8060 => x"00000016", -- pedding 
        8061 => x"00000016", -- pedding 
        8062 => x"00000016", -- pedding 
        8063 => x"00000016", -- pedding 
        8064 => x"00000016", -- pedding 
        8065 => x"00000016", -- pedding 
        8066 => x"00000016", -- pedding 
        8067 => x"00000016", -- pedding 
        8068 => x"00000016", -- pedding 
        8069 => x"00000016", -- pedding 
        8070 => x"00000016", -- pedding 
        8071 => x"00000016", -- pedding 
        8072 => x"00000016", -- pedding 
        8073 => x"00000016", -- pedding 
        8074 => x"00000016", -- pedding 
        8075 => x"00000016", -- pedding 
        8076 => x"00000016", -- pedding 
        8077 => x"00000016", -- pedding 
        8078 => x"00000016", -- pedding 
        8079 => x"00000016", -- pedding 
        8080 => x"00000016", -- pedding 
        8081 => x"00000016", -- pedding 
        8082 => x"00000016", -- pedding 
        8083 => x"00000016", -- pedding 
        8084 => x"00000016", -- pedding 
        8085 => x"00000016", -- pedding 
        8086 => x"00000016", -- pedding 
        8087 => x"00000016", -- pedding 
        8088 => x"00000016", -- pedding 
        8089 => x"00000016", -- pedding 
        8090 => x"00000016", -- pedding 
        8091 => x"00000016", -- pedding 
        8092 => x"00000016", -- pedding 
        8093 => x"00000016", -- pedding 
        8094 => x"00000016", -- pedding 
        8095 => x"00000016", -- pedding 
        8096 => x"00000016", -- pedding 
        8097 => x"00000016", -- pedding 
        8098 => x"00000016", -- pedding 
        8099 => x"00000016", -- pedding 
        8100 => x"00000016", -- pedding 
        8101 => x"00000016", -- pedding 
        8102 => x"00000016", -- pedding 
        8103 => x"00000016", -- pedding 
        8104 => x"00000016", -- pedding 
        8105 => x"00000016", -- pedding 
        8106 => x"00000016", -- pedding 
        8107 => x"00000016", -- pedding 
        8108 => x"00000016", -- pedding 
        8109 => x"00000016", -- pedding 
        8110 => x"00000016", -- pedding 
        8111 => x"00000016", -- pedding 
        8112 => x"00000016", -- pedding 
        8113 => x"00000016", -- pedding 
        8114 => x"00000016", -- pedding 
        8115 => x"00000016", -- pedding 
        8116 => x"00000016", -- pedding 
        8117 => x"00000016", -- pedding 
        8118 => x"00000016", -- pedding 
        8119 => x"00000016", -- pedding 
        8120 => x"00000016", -- pedding 
        8121 => x"00000016", -- pedding 
        8122 => x"00000016", -- pedding 
        8123 => x"00000016", -- pedding 
        8124 => x"00000016", -- pedding 
        8125 => x"00000016", -- pedding 
        8126 => x"00000016", -- pedding 
        8127 => x"00000016", -- pedding 
        8128 => x"00000016", -- pedding 
        8129 => x"00000016", -- pedding 
        8130 => x"00000016", -- pedding 
        8131 => x"00000016", -- pedding 
        8132 => x"00000016", -- pedding 
        8133 => x"00000016", -- pedding 
        8134 => x"00000016", -- pedding 
        8135 => x"00000016", -- pedding 
        8136 => x"00000016", -- pedding 
        8137 => x"00000016", -- pedding 
        8138 => x"00000016", -- pedding 
        8139 => x"00000016", -- pedding 
        8140 => x"00000016", -- pedding 
        8141 => x"00000016", -- pedding 
        8142 => x"00000016", -- pedding 
        8143 => x"00000016", -- pedding 
        8144 => x"00000016", -- pedding 
        8145 => x"00000016", -- pedding 
        8146 => x"00000016", -- pedding 
        8147 => x"00000016", -- pedding 
        8148 => x"00000016", -- pedding 
        8149 => x"00000016", -- pedding 
        8150 => x"00000016", -- pedding 
        8151 => x"00000016", -- pedding 
        8152 => x"00000016", -- pedding 
        8153 => x"00000016", -- pedding 
        8154 => x"00000016", -- pedding 
        8155 => x"00000016", -- pedding 
        8156 => x"00000016", -- pedding 
        8157 => x"00000016", -- pedding 
        8158 => x"00000016", -- pedding 
        8159 => x"00000016", -- pedding 
        8160 => x"00000016", -- pedding 
        8161 => x"00000016", -- pedding 
        8162 => x"00000016", -- pedding 
        8163 => x"00000016", -- pedding 
        8164 => x"00000016", -- pedding 
        8165 => x"00000016", -- pedding 
        8166 => x"00000016", -- pedding 
        8167 => x"00000016", -- pedding 
        8168 => x"00000016", -- pedding 
        8169 => x"00000016", -- pedding 
        8170 => x"00000016", -- pedding 
        8171 => x"00000016", -- pedding 
        8172 => x"00000016", -- pedding 
        8173 => x"00000016", -- pedding 
        8174 => x"00000016", -- pedding 
        8175 => x"00000016", -- pedding 
        8176 => x"00000016", -- pedding 
        8177 => x"00000016", -- pedding 
        8178 => x"00000016", -- pedding 
        8179 => x"00000016", -- pedding 
        8180 => x"00000016", -- pedding 
        8181 => x"00000016", -- pedding 
        8182 => x"00000016", -- pedding 
        8183 => x"00000016", -- pedding 
        8184 => x"00000016", -- pedding 
        8185 => x"00000016", -- pedding 
        8186 => x"00000016", -- pedding 
        8187 => x"00000016", -- pedding 
        8188 => x"00000016", -- pedding 
        8189 => x"00000016", -- pedding 
        8190 => x"00000016", -- pedding 
        8191 => x"00000016", -- pedding


others => x"00000000"
	);


begin

	process(i_clk)
	begin
		if rising_edge(i_clk) then
			-- memory write --
			if i_we = '1' then
				mem(to_integer(unsigned(i_w_addr))) <= i_data;
			end if;
			-- memory read --
			o_data <= mem(to_integer(unsigned(i_r_addr)));

		end if;
	end process;

end architecture arch;
