library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity ram is
	generic
	(
		DATA_WIDTH : natural := 32;		    -- 4 byte one line of memory
		ADDR_WIDTH : natural := 13			    -- 24576 bytes size of memory
	);

	port(
		i_clk    : in  std_logic;
		i_r_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		i_data   : in  std_logic_vector(DATA_WIDTH-1 downto 0);
		i_we     : in  std_logic;
		i_w_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		o_data   : out std_logic_vector(DATA_WIDTH-1 downto 0)
	);
end entity ram;

architecture arch of ram is

	type ram_t is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(DATA_WIDTH-1 downto 0);


-- GENERATED BY BC_MEM_PACKER

-- DATE: Thu May 18 16:01:02 2017

	signal mem : ram_t := (

--			***** COLOR PALLETE *****

		-- fellas
		0 =>	x"00000000",
		1 =>	x"00A8D8FC",
		2 =>	x"00000000",
		3 =>	x"00EC3820",
		4 =>	x"0000A800",
		5 =>	x"00FCFCFC",
		6 =>	x"00747474",
		7 =>	x"00C0C0C0",
--      Link colors

        8 =>      x"00303030",
        9 =>      x"000CCB83",
        10 =>     x"002C98D8",
        11 =>     x"00004B7B",
        12 =>     x"00FFD9D9",
        13 =>     x"00003299",
        14 =>     x"00B1DFF8",
        15 =>     x"00FFFFFF",
        16 =>     x"008E0018",
        17 =>     x"00FF898E",
        18 =>     x"00000000",
        19 =>     x"00006E8A",
        20 =>     x"00002E55",
        21 =>     x"00CBC74D",
        22 =>     x"00E32F47",
        23 =>     x"00173B00",
        24 =>     x"00007A3E",
        25 =>     x"007ED14A",
        26 =>     x"0000311D",
        27 =>     x"0000675B",
        28 =>     x"000AB4B9",
        29 =>     x"00003D00",
        30 =>     x"00008200",
        31 =>     x"003FD65B",
        32 =>     x"00656565",
        33 =>     x"00B9B9B9",
        34 =>     x"00AFAFAF",

        

-- 		vatrie colors

  35=>    x"00000000",
  36=>    x"000038f8",
  37=>    x"00abe3ff",
  38=>    x"00ffffff",
		-- map colors

40=> x"00bc0000",
41=> x"00000000",
42=> x"0044a0fc",
43=> x"00d8e800",

-- majmun1 colors
  44=>    x"00000000",
  45=>    x"000013ab",
  46=>    x"00b0d0F0",
  47=>    x"00ffffff",
-- majmun2 colors
  --48=>    x"00000000",
  48=>    x"00000000",
  49=>    x"000013ab",
  50=>    x"00b0d0F0",
  51=>    x"00ffffff",

--mario colors
  52=>    x"00000000",
  --52=>    x"00ffffff",
  53=>    x"000000ff",
  54=>    x"009cd0ea",
  55=>    x"00db0000",

--princeza colors

56=>    x"00000000",
57=>    x"004e4e76",
58=>    x"00bbe4f9",
59=>    x"00ff00ff",

		60 => x"00000000",
		61 => x"00000203",
		62 => x"000000ff",



	63 =>	x"003199FF", -- Unused

            --  ADDED SPRITES HERE
          -- RUPEE SPRITE
		64 => x"0202020F",
		65 => x"3C020202",
		66 => x"02020202",
		67 => x"02020202",
		68 => x"02020F0F",
		69 => x"3C3C0202",
		70 => x"02020202",
		71 => x"02020202",
		72 => x"020F0F0F",
		73 => x"3C3C3C02",
		74 => x"02020202",
		75 => x"02020202",
		76 => x"0F3C0F3C",
		77 => x"023C023C",
		78 => x"02020202",
		79 => x"02020202",
		80 => x"0F0F3C3C",
		81 => x"3C023C3C",
		82 => x"02020202",
		83 => x"02020202",
		84 => x"0F0F3C3C",
		85 => x"3C023C3C",
		86 => x"02020202",
		87 => x"02020202",
		88 => x"0F0F3C3C",
		89 => x"3C023C3C",
		90 => x"02020202",
		91 => x"02020202",
		92 => x"0F0F3C3C",
		93 => x"3C023C3C",
		94 => x"02020202",
		95 => x"02020202",
		96 => x"0F0F3C3C",
		97 => x"3C023C3C",
		98 => x"02020202",
		99 => x"02020202",
		100 => x"0F0F3C3C",
		101 => x"3C023C3C",
		102 => x"02020202",
		103 => x"02020202",
		104 => x"0F0F3C3C",
		105 => x"3C023C3C",
		106 => x"02020202",
		107 => x"02020202",
		108 => x"0F3C0F3C",
		109 => x"3C023C3C",
		110 => x"02020202",
		111 => x"02020202",
		112 => x"3C3C3C0F",
		113 => x"023C023C",
		114 => x"02020202",
		115 => x"02020202",
		116 => x"023C3C3C",
		117 => x"3C3C3C02",
		118 => x"02020202",
		119 => x"02020202",
		120 => x"02023C3C",
		121 => x"3C3C0202",
		122 => x"02020202",
		123 => x"02020202",
		124 => x"0202023C",
		125 => x"3C020202",
		126 => x"02020202",
		127 => x"02020202",

          -- BOMB SPRITE
		128 => x"02020202",
		129 => x"020F0202",
		130 => x"02020202",
		131 => x"02020202",
		132 => x"02020202",
		133 => x"020F0202",
		134 => x"02020202",
		135 => x"02020202",
		136 => x"02020202",
		137 => x"02020F02",
		138 => x"02020202",
		139 => x"02020202",
		140 => x"02020202",
		141 => x"0202020F",
		142 => x"02020202",
		143 => x"02020202",
		144 => x"02020202",
		145 => x"0202020F",
		146 => x"02020202",
		147 => x"02020202",
		148 => x"02020202",
		149 => x"02020F02",
		150 => x"02020202",
		151 => x"02020202",
		152 => x"02020D0D",
		153 => x"0D0D0202",
		154 => x"02020202",
		155 => x"02020202",
		156 => x"020D2E2E",
		157 => x"0D0D0D02",
		158 => x"02020202",
		159 => x"02020202",
		160 => x"0D2E0F2E",
		161 => x"0D0D0D0D",
		162 => x"02020202",
		163 => x"02020202",
		164 => x"0D2E2E0D",
		165 => x"0D0D0D0D",
		166 => x"02020202",
		167 => x"02020202",
		168 => x"0D0D0D0D",
		169 => x"0D0D0D0D",
		170 => x"02020202",
		171 => x"02020202",
		172 => x"0D0D0D0D",
		173 => x"0D0D0D0D",
		174 => x"02020202",
		175 => x"02020202",
		176 => x"020D0D0D",
		177 => x"0D0D0D02",
		178 => x"02020202",
		179 => x"02020202",
		180 => x"02020D0D",
		181 => x"0D0D0202",
		182 => x"02020202",
		183 => x"02020202",
		184 => x"02020202",
		185 => x"02020202",
		186 => x"02020202",
		187 => x"02020202",
		188 => x"02020202",
		189 => x"02020202",
		190 => x"02020202",
		191 => x"02020202",
		
		--Trambolina
		  192 => x"29292929",		-- colors: 41, 41, 41, 41
        193 => x"29292929",		-- colors: 41, 41, 41, 41
        194 => x"29292929",		-- colors: 41, 41, 41, 41
        195 => x"29292929",		-- colors: 41, 41, 41, 41
        196 => x"29292929",		-- colors: 41, 41, 41, 41
        197 => x"29292929",		-- colors: 41, 41, 41, 41
        198 => x"29292929",		-- colors: 41, 41, 41, 41
        199 => x"29292929",		-- colors: 41, 41, 41, 41
        200 => x"29292929",		-- colors: 41, 41, 41, 41
        201 => x"24242424",		-- colors: 41, 41, 41, 41
        202 => x"24242424",		-- colors: 41, 41, 41, 41
        203 => x"29292929",		-- colors: 41, 41, 41, 41
        204 => x"29292929",		-- colors: 41, 41, 41, 41
        205 => x"24242424",		-- colors: 41, 41, 41, 41
        206 => x"24242424",		-- colors: 41, 41, 41, 41
        207 => x"29292929",		-- colors: 41, 41, 41, 41
        208 => x"28282828",		-- colors: 41, 41, 41, 41
        209 => x"28282828",		-- colors: 41, 41, 41, 41
        210 => x"28282828",		-- colors: 41, 41, 41, 41
        211 => x"28282828",		-- colors: 41, 41, 41, 41
        212 => x"28282828",		-- colors: 41, 41, 41, 41
        213 => x"28282828",		-- colors: 41, 41, 41, 41
        214 => x"28282828",		-- colors: 41, 41, 41, 41
        215 => x"28282828",		-- colors: 41, 41, 41, 41
        216 => x"28282828",		-- colors: 41, 41, 41, 41
        217 => x"28282828",		-- colors: 41, 41, 41, 41
        218 => x"28282828",		-- colors: 41, 41, 41, 41
        219 => x"28282828",		-- colors: 41, 41, 41, 41
        220 => x"28282828",		-- colors: 41, 41, 41, 41
        221 => x"28282828",		-- colors: 41, 41, 41, 41
        222 => x"28282828",		-- colors: 41, 41, 41, 41
        223 => x"28282828",		-- colors: 41, 41, 41, 41
        224 => x"28282828",		-- colors: 40, 40, 40, 40
        225 => x"28282828",		-- colors: 40, 40, 40, 40
        226 => x"28282828",		-- colors: 40, 40, 40, 40
        227 => x"28282828",		-- colors: 40, 40, 40, 40
        228 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        229 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        230 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        231 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        232 => x"28282929",		-- colors: 40, 40, 41, 41
        233 => x"29292828",		-- colors: 41, 41, 40, 40
        234 => x"28282929",		-- colors: 40, 40, 41, 41
        235 => x"29292828",		-- colors: 41, 41, 40, 40
        236 => x"28292929",		-- colors: 40, 41, 41, 41
        237 => x"29292928",		-- colors: 41, 41, 41, 40
        238 => x"28292929",		-- colors: 40, 41, 41, 41
        239 => x"29292928",		-- colors: 41, 41, 41, 40
        240 => x"28292929",		-- colors: 40, 41, 41, 41
        241 => x"29292928",		-- colors: 41, 41, 41, 40
        242 => x"28292929",		-- colors: 40, 41, 41, 41
        243 => x"29292928",		-- colors: 41, 41, 41, 40
        244 => x"28282929",		-- colors: 40, 40, 41, 41
        245 => x"29292828",		-- colors: 41, 41, 40, 40
        246 => x"28282929",		-- colors: 40, 40, 41, 41
        247 => x"29292828",		-- colors: 41, 41, 40, 40
        248 => x"28282828",		-- colors: 40, 40, 40, 40
        249 => x"28282828",		-- colors: 40, 40, 40, 40
        250 => x"28282828",		-- colors: 40, 40, 40, 40
        251 => x"28282828",		-- colors: 40, 40, 40, 40
        252 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        253 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        254 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        
        

--			***** 16x16 IMAGES *****
--			OVERWORLD SPRITES
  --  sprite 0
        255 => x"28282828",		-- colors: 40, 40, 40, 40
        256 => x"28282828",		-- colors: 40, 40, 40, 40
        257 => x"28282828",		-- colors: 40, 40, 40, 40
        258 => x"28282828",		-- colors: 40, 40, 40, 40
        259 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        260 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        261 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        262 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        263 => x"28282929",		-- colors: 40, 40, 41, 41
        264 => x"29292828",		-- colors: 41, 41, 40, 40
        265 => x"28282929",		-- colors: 40, 40, 41, 41
        266 => x"29292828",		-- colors: 41, 41, 40, 40
        267 => x"28292929",		-- colors: 40, 41, 41, 41
        268 => x"29292928",		-- colors: 41, 41, 41, 40
        269 => x"28292929",		-- colors: 40, 41, 41, 41
        270 => x"29292928",		-- colors: 41, 41, 41, 40
        271 => x"28292929",		-- colors: 40, 41, 41, 41
        272 => x"29292928",		-- colors: 41, 41, 41, 40
        273 => x"28292929",		-- colors: 40, 41, 41, 41
        274 => x"29292928",		-- colors: 41, 41, 41, 40
        275 => x"28282929",		-- colors: 40, 40, 41, 41
        276 => x"29292828",		-- colors: 41, 41, 40, 40
        277 => x"28282929",		-- colors: 40, 40, 41, 41
        278 => x"29292828",		-- colors: 41, 41, 40, 40
        279 => x"28282828",		-- colors: 40, 40, 40, 40
        280 => x"28282828",		-- colors: 40, 40, 40, 40
        281 => x"28282828",		-- colors: 40, 40, 40, 40
        282 => x"28282828",		-- colors: 40, 40, 40, 40
        283 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        284 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        285 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        286 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        287 => x"29292929",		-- colors: 41, 41, 41, 41
        288 => x"29292929",		-- colors: 41, 41, 41, 41
        289 => x"29292929",		-- colors: 41, 41, 41, 41
        290 => x"29292929",		-- colors: 41, 41, 41, 41
        291 => x"29292929",		-- colors: 41, 41, 41, 41
        292 => x"29292929",		-- colors: 41, 41, 41, 41
        293 => x"29292929",		-- colors: 41, 41, 41, 41
        294 => x"29292929",		-- colors: 41, 41, 41, 41
        295 => x"29292929",		-- colors: 41, 41, 41, 41
        296 => x"29292929",		-- colors: 41, 41, 41, 41
        297 => x"29292929",		-- colors: 41, 41, 41, 41
        298 => x"29292929",		-- colors: 41, 41, 41, 41
        299 => x"29292929",		-- colors: 41, 41, 41, 41
        300 => x"29292929",		-- colors: 41, 41, 41, 41
        301 => x"29292929",		-- colors: 41, 41, 41, 41
        302 => x"29292929",		-- colors: 41, 41, 41, 41
        303 => x"29292929",		-- colors: 41, 41, 41, 41
        304 => x"29292929",		-- colors: 41, 41, 41, 41
        305 => x"29292929",		-- colors: 41, 41, 41, 41
        306 => x"29292929",		-- colors: 41, 41, 41, 41
        307 => x"29292929",		-- colors: 41, 41, 41, 41
        308 => x"29292929",		-- colors: 41, 41, 41, 41
        309 => x"29292929",		-- colors: 41, 41, 41, 41
        310 => x"29292929",		-- colors: 41, 41, 41, 41
        311 => x"29292929",		-- colors: 41, 41, 41, 41
        312 => x"29292929",		-- colors: 41, 41, 41, 41
        313 => x"29292929",		-- colors: 41, 41, 41, 41
        314 => x"29292929",		-- colors: 41, 41, 41, 41
        315 => x"29292929",		-- colors: 41, 41, 41, 41
        316 => x"29292929",		-- colors: 41, 41, 41, 41
        317 => x"29292929",		-- colors: 41, 41, 41, 41
        318 => x"29292929",		-- colors: 41, 41, 41, 41

                --  sprite 1
        319 => x"29292929",		-- colors: 41, 41, 41, 41
        320 => x"29292929",		-- colors: 41, 41, 41, 41
        321 => x"29292929",		-- colors: 41, 41, 41, 41
        322 => x"29292929",		-- colors: 41, 41, 41, 41
        323 => x"29292929",		-- colors: 41, 41, 41, 41
        324 => x"29292929",		-- colors: 41, 41, 41, 41
        325 => x"29292929",		-- colors: 41, 41, 41, 41
        326 => x"29292929",		-- colors: 41, 41, 41, 41
        327 => x"29292929",		-- colors: 41, 41, 41, 41
        328 => x"29292929",		-- colors: 41, 41, 41, 41
        329 => x"29292929",		-- colors: 41, 41, 41, 41
        330 => x"29292929",		-- colors: 41, 41, 41, 41
        331 => x"29292929",		-- colors: 41, 41, 41, 41
        332 => x"29292929",		-- colors: 41, 41, 41, 41
        333 => x"29292929",		-- colors: 41, 41, 41, 41
        334 => x"29292929",		-- colors: 41, 41, 41, 41
        335 => x"29292929",		-- colors: 41, 41, 41, 41
        336 => x"29292929",		-- colors: 41, 41, 41, 41
        337 => x"29292929",		-- colors: 41, 41, 41, 41
        338 => x"29292929",		-- colors: 41, 41, 41, 41
        339 => x"29292929",		-- colors: 41, 41, 41, 41
        340 => x"29292929",		-- colors: 41, 41, 41, 41
        341 => x"29292929",		-- colors: 41, 41, 41, 41
        342 => x"29292929",		-- colors: 41, 41, 41, 41
        343 => x"29292929",		-- colors: 41, 41, 41, 41
        344 => x"29292929",		-- colors: 41, 41, 41, 41
        345 => x"29292929",		-- colors: 41, 41, 41, 41
        346 => x"29292929",		-- colors: 41, 41, 41, 41
        347 => x"29292929",		-- colors: 41, 41, 41, 41
        348 => x"29292929",		-- colors: 41, 41, 41, 41
        349 => x"29292929",		-- colors: 41, 41, 41, 41
        350 => x"29292929",		-- colors: 41, 41, 41, 41
        351 => x"28282828",		-- colors: 40, 40, 40, 40
        352 => x"28282828",		-- colors: 40, 40, 40, 40
        353 => x"28282828",		-- colors: 40, 40, 40, 40
        354 => x"28282828",		-- colors: 40, 40, 40, 40
        355 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        356 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        357 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        358 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        359 => x"28282929",		-- colors: 40, 40, 41, 41
        360 => x"29292828",		-- colors: 41, 41, 40, 40
        361 => x"28282929",		-- colors: 40, 40, 41, 41
        362 => x"29292828",		-- colors: 41, 41, 40, 40
        363 => x"28292929",		-- colors: 40, 41, 41, 41
        364 => x"29292928",		-- colors: 41, 41, 41, 40
        365 => x"28292929",		-- colors: 40, 41, 41, 41
        366 => x"29292928",		-- colors: 41, 41, 41, 40
        367 => x"28292929",		-- colors: 40, 41, 41, 41
        368 => x"29292928",		-- colors: 41, 41, 41, 40
        369 => x"28292929",		-- colors: 40, 41, 41, 41
        370 => x"29292928",		-- colors: 41, 41, 41, 40
        371 => x"28282929",		-- colors: 40, 40, 41, 41
        372 => x"29292828",		-- colors: 41, 41, 40, 40
        373 => x"28282929",		-- colors: 40, 40, 41, 41
        374 => x"29292828",		-- colors: 41, 41, 40, 40
        375 => x"28282828",		-- colors: 40, 40, 40, 40
        376 => x"28282828",		-- colors: 40, 40, 40, 40
        377 => x"28282828",		-- colors: 40, 40, 40, 40
        378 => x"28282828",		-- colors: 40, 40, 40, 40
        379 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        380 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        381 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        382 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43

                --  sprite 2
        383 => x"29292929",		-- colors: 41, 41, 41, 41
        384 => x"29292929",		-- colors: 41, 41, 41, 41
        385 => x"2A292929",		-- colors: 42, 41, 41, 41
        386 => x"2929292A",		-- colors: 41, 41, 41, 42
        387 => x"29292929",		-- colors: 41, 41, 41, 41
        388 => x"29292929",		-- colors: 41, 41, 41, 41
        389 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
        390 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
        391 => x"29292929",		-- colors: 41, 41, 41, 41
        392 => x"29292929",		-- colors: 41, 41, 41, 41
        393 => x"2A292929",		-- colors: 42, 41, 41, 41
        394 => x"2929292A",		-- colors: 41, 41, 41, 42
        395 => x"29292929",		-- colors: 41, 41, 41, 41
        396 => x"29292929",		-- colors: 41, 41, 41, 41
        397 => x"2A292929",		-- colors: 42, 41, 41, 41
        398 => x"2929292A",		-- colors: 41, 41, 41, 42
        399 => x"29292929",		-- colors: 41, 41, 41, 41
        400 => x"29292929",		-- colors: 41, 41, 41, 41
        401 => x"2A292929",		-- colors: 42, 41, 41, 41
        402 => x"2929292A",		-- colors: 41, 41, 41, 42
        403 => x"29292929",		-- colors: 41, 41, 41, 41
        404 => x"29292929",		-- colors: 41, 41, 41, 41
        405 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
        406 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
        407 => x"29292929",		-- colors: 41, 41, 41, 41
        408 => x"29292929",		-- colors: 41, 41, 41, 41
        409 => x"2A292929",		-- colors: 42, 41, 41, 41
        410 => x"2929292A",		-- colors: 41, 41, 41, 42
        411 => x"29292929",		-- colors: 41, 41, 41, 41
        412 => x"29292929",		-- colors: 41, 41, 41, 41
        413 => x"2A292929",		-- colors: 42, 41, 41, 41
        414 => x"2929292A",		-- colors: 41, 41, 41, 42
        415 => x"28282828",		-- colors: 40, 40, 40, 40
        416 => x"28282828",		-- colors: 40, 40, 40, 40
        417 => x"28282828",		-- colors: 40, 40, 40, 40
        418 => x"28282828",		-- colors: 40, 40, 40, 40
        419 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        420 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        421 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        422 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        423 => x"28282929",		-- colors: 40, 40, 41, 41
        424 => x"29292828",		-- colors: 41, 41, 40, 40
        425 => x"28282929",		-- colors: 40, 40, 41, 41
        426 => x"29292828",		-- colors: 41, 41, 40, 40
        427 => x"28292929",		-- colors: 40, 41, 41, 41
        428 => x"29292928",		-- colors: 41, 41, 41, 40
        429 => x"28292929",		-- colors: 40, 41, 41, 41
        430 => x"29292928",		-- colors: 41, 41, 41, 40
        431 => x"28292929",		-- colors: 40, 41, 41, 41
        432 => x"29292928",		-- colors: 41, 41, 41, 40
        433 => x"28292929",		-- colors: 40, 41, 41, 41
        434 => x"29292928",		-- colors: 41, 41, 41, 40
        435 => x"28282929",		-- colors: 40, 40, 41, 41
        436 => x"29292828",		-- colors: 41, 41, 40, 40
        437 => x"28282929",		-- colors: 40, 40, 41, 41
        438 => x"29292828",		-- colors: 41, 41, 40, 40
        439 => x"28282828",		-- colors: 40, 40, 40, 40
        440 => x"28282828",		-- colors: 40, 40, 40, 40
        441 => x"28282828",		-- colors: 40, 40, 40, 40
        442 => x"28282828",		-- colors: 40, 40, 40, 40
        443 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        444 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        445 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        446 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43

                --  sprite 3
        447 => x"2A292929",		-- colors: 42, 41, 41, 41
        448 => x"2929292A",		-- colors: 41, 41, 41, 42
        449 => x"29292929",		-- colors: 41, 41, 41, 41
        450 => x"29292929",		-- colors: 41, 41, 41, 41
        451 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
        452 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
        453 => x"29292929",		-- colors: 41, 41, 41, 41
        454 => x"29292929",		-- colors: 41, 41, 41, 41
        455 => x"2A292929",		-- colors: 42, 41, 41, 41
        456 => x"2929292A",		-- colors: 41, 41, 41, 42
        457 => x"29292929",		-- colors: 41, 41, 41, 41
        458 => x"29292929",		-- colors: 41, 41, 41, 41
        459 => x"2A292929",		-- colors: 42, 41, 41, 41
        460 => x"2929292A",		-- colors: 41, 41, 41, 42
        461 => x"29292929",		-- colors: 41, 41, 41, 41
        462 => x"29292929",		-- colors: 41, 41, 41, 41
        463 => x"2A292929",		-- colors: 42, 41, 41, 41
        464 => x"2929292A",		-- colors: 41, 41, 41, 42
        465 => x"29292929",		-- colors: 41, 41, 41, 41
        466 => x"29292929",		-- colors: 41, 41, 41, 41
        467 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
        468 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
        469 => x"29292929",		-- colors: 41, 41, 41, 41
        470 => x"29292929",		-- colors: 41, 41, 41, 41
        471 => x"2A292929",		-- colors: 42, 41, 41, 41
        472 => x"2929292A",		-- colors: 41, 41, 41, 42
        473 => x"29292929",		-- colors: 41, 41, 41, 41
        474 => x"29292929",		-- colors: 41, 41, 41, 41
        475 => x"2A292929",		-- colors: 42, 41, 41, 41
        476 => x"2929292A",		-- colors: 41, 41, 41, 42
        477 => x"29292929",		-- colors: 41, 41, 41, 41
        478 => x"29292929",		-- colors: 41, 41, 41, 41
        479 => x"28282828",		-- colors: 40, 40, 40, 40
        480 => x"28282828",		-- colors: 40, 40, 40, 40
        481 => x"28282828",		-- colors: 40, 40, 40, 40
        482 => x"28282828",		-- colors: 40, 40, 40, 40
        483 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        484 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        485 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        486 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        487 => x"28282929",		-- colors: 40, 40, 41, 41
        488 => x"29292828",		-- colors: 41, 41, 40, 40
        489 => x"28282929",		-- colors: 40, 40, 41, 41
        490 => x"29292828",		-- colors: 41, 41, 40, 40
        491 => x"28292929",		-- colors: 40, 41, 41, 41
        492 => x"29292928",		-- colors: 41, 41, 41, 40
        493 => x"28292929",		-- colors: 40, 41, 41, 41
        494 => x"29292928",		-- colors: 41, 41, 41, 40
        495 => x"28292929",		-- colors: 40, 41, 41, 41
        496 => x"29292928",		-- colors: 41, 41, 41, 40
        497 => x"28292929",		-- colors: 40, 41, 41, 41
        498 => x"29292928",		-- colors: 41, 41, 41, 40
        499 => x"28282929",		-- colors: 40, 40, 41, 41
        500 => x"29292828",		-- colors: 41, 41, 40, 40
        501 => x"28282929",		-- colors: 40, 40, 41, 41
        502 => x"29292828",		-- colors: 41, 41, 40, 40
        503 => x"28282828",		-- colors: 40, 40, 40, 40
        504 => x"28282828",		-- colors: 40, 40, 40, 40
        505 => x"28282828",		-- colors: 40, 40, 40, 40
        506 => x"28282828",		-- colors: 40, 40, 40, 40
        507 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        508 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        509 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        510 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43

                --  sprite 4
        511 => x"2A292929",		-- colors: 42, 41, 41, 41
        512 => x"2929292A",		-- colors: 41, 41, 41, 42
        513 => x"29292929",		-- colors: 41, 41, 41, 41
        514 => x"29292929",		-- colors: 41, 41, 41, 41
        515 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
        516 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
        517 => x"29292929",		-- colors: 41, 41, 41, 41
        518 => x"29292929",		-- colors: 41, 41, 41, 41
        519 => x"2A292929",		-- colors: 42, 41, 41, 41
        520 => x"2929292A",		-- colors: 41, 41, 41, 42
        521 => x"29292929",		-- colors: 41, 41, 41, 41
        522 => x"29292929",		-- colors: 41, 41, 41, 41
        523 => x"2A292929",		-- colors: 42, 41, 41, 41
        524 => x"2929292A",		-- colors: 41, 41, 41, 42
        525 => x"29292929",		-- colors: 41, 41, 41, 41
        526 => x"29292929",		-- colors: 41, 41, 41, 41
        527 => x"2A292929",		-- colors: 42, 41, 41, 41
        528 => x"2929292A",		-- colors: 41, 41, 41, 42
        529 => x"29292929",		-- colors: 41, 41, 41, 41
        530 => x"29292929",		-- colors: 41, 41, 41, 41
        531 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
        532 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
        533 => x"29292929",		-- colors: 41, 41, 41, 41
        534 => x"29292929",		-- colors: 41, 41, 41, 41
        535 => x"2A292929",		-- colors: 42, 41, 41, 41
        536 => x"2929292A",		-- colors: 41, 41, 41, 42
        537 => x"29292929",		-- colors: 41, 41, 41, 41
        538 => x"29292929",		-- colors: 41, 41, 41, 41
        539 => x"2A292929",		-- colors: 42, 41, 41, 41
        540 => x"2929292A",		-- colors: 41, 41, 41, 42
        541 => x"29292929",		-- colors: 41, 41, 41, 41
        542 => x"29292929",		-- colors: 41, 41, 41, 41
        543 => x"2A292929",		-- colors: 42, 41, 41, 41
        544 => x"2929292A",		-- colors: 41, 41, 41, 42
        545 => x"29292929",		-- colors: 41, 41, 41, 41
        546 => x"29292929",		-- colors: 41, 41, 41, 41
        547 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
        548 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
        549 => x"29292929",		-- colors: 41, 41, 41, 41
        550 => x"29292929",		-- colors: 41, 41, 41, 41
        551 => x"2A292929",		-- colors: 42, 41, 41, 41
        552 => x"2929292A",		-- colors: 41, 41, 41, 42
        553 => x"29292929",		-- colors: 41, 41, 41, 41
        554 => x"29292929",		-- colors: 41, 41, 41, 41
        555 => x"2A292929",		-- colors: 42, 41, 41, 41
        556 => x"2929292A",		-- colors: 41, 41, 41, 42
        557 => x"29292929",		-- colors: 41, 41, 41, 41
        558 => x"29292929",		-- colors: 41, 41, 41, 41
        559 => x"2A292929",		-- colors: 42, 41, 41, 41
        560 => x"2929292A",		-- colors: 41, 41, 41, 42
        561 => x"29292929",		-- colors: 41, 41, 41, 41
        562 => x"29292929",		-- colors: 41, 41, 41, 41
        563 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
        564 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
        565 => x"29292929",		-- colors: 41, 41, 41, 41
        566 => x"29292929",		-- colors: 41, 41, 41, 41
        567 => x"2A292929",		-- colors: 42, 41, 41, 41
        568 => x"2929292A",		-- colors: 41, 41, 41, 42
        569 => x"29292929",		-- colors: 41, 41, 41, 41
        570 => x"29292929",		-- colors: 41, 41, 41, 41
        571 => x"2A292929",		-- colors: 42, 41, 41, 41
        572 => x"2929292A",		-- colors: 41, 41, 41, 42
        573 => x"29292929",		-- colors: 41, 41, 41, 41
        574 => x"29292929",		-- colors: 41, 41, 41, 41

                --  sprite 5
        575 => x"29292929",		-- colors: 41, 41, 41, 41
        576 => x"29292929",		-- colors: 41, 41, 41, 41
        577 => x"2A292929",		-- colors: 42, 41, 41, 41
        578 => x"2929292A",		-- colors: 41, 41, 41, 42
        579 => x"29292929",		-- colors: 41, 41, 41, 41
        580 => x"29292929",		-- colors: 41, 41, 41, 41
        581 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
        582 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
        583 => x"29292929",		-- colors: 41, 41, 41, 41
        584 => x"29292929",		-- colors: 41, 41, 41, 41
        585 => x"2A292929",		-- colors: 42, 41, 41, 41
        586 => x"2929292A",		-- colors: 41, 41, 41, 42
        587 => x"29292929",		-- colors: 41, 41, 41, 41
        588 => x"29292929",		-- colors: 41, 41, 41, 41
        589 => x"2A292929",		-- colors: 42, 41, 41, 41
        590 => x"2929292A",		-- colors: 41, 41, 41, 42
        591 => x"29292929",		-- colors: 41, 41, 41, 41
        592 => x"29292929",		-- colors: 41, 41, 41, 41
        593 => x"2A292929",		-- colors: 42, 41, 41, 41
        594 => x"2929292A",		-- colors: 41, 41, 41, 42
        595 => x"29292929",		-- colors: 41, 41, 41, 41
        596 => x"29292929",		-- colors: 41, 41, 41, 41
        597 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
        598 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
        599 => x"29292929",		-- colors: 41, 41, 41, 41
        600 => x"29292929",		-- colors: 41, 41, 41, 41
        601 => x"2A292929",		-- colors: 42, 41, 41, 41
        602 => x"2929292A",		-- colors: 41, 41, 41, 42
        603 => x"29292929",		-- colors: 41, 41, 41, 41
        604 => x"29292929",		-- colors: 41, 41, 41, 41
        605 => x"2A292929",		-- colors: 42, 41, 41, 41
        606 => x"2929292A",		-- colors: 41, 41, 41, 42
        607 => x"29292929",		-- colors: 41, 41, 41, 41
        608 => x"29292929",		-- colors: 41, 41, 41, 41
        609 => x"2A292929",		-- colors: 42, 41, 41, 41
        610 => x"2929292A",		-- colors: 41, 41, 41, 42
        611 => x"29292929",		-- colors: 41, 41, 41, 41
        612 => x"29292929",		-- colors: 41, 41, 41, 41
        613 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
        614 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
        615 => x"29292929",		-- colors: 41, 41, 41, 41
        616 => x"29292929",		-- colors: 41, 41, 41, 41
        617 => x"2A292929",		-- colors: 42, 41, 41, 41
        618 => x"2929292A",		-- colors: 41, 41, 41, 42
        619 => x"29292929",		-- colors: 41, 41, 41, 41
        620 => x"29292929",		-- colors: 41, 41, 41, 41
        621 => x"2A292929",		-- colors: 42, 41, 41, 41
        622 => x"2929292A",		-- colors: 41, 41, 41, 42
        623 => x"29292929",		-- colors: 41, 41, 41, 41
        624 => x"29292929",		-- colors: 41, 41, 41, 41
        625 => x"2A292929",		-- colors: 42, 41, 41, 41
        626 => x"2929292A",		-- colors: 41, 41, 41, 42
        627 => x"29292929",		-- colors: 41, 41, 41, 41
        628 => x"29292929",		-- colors: 41, 41, 41, 41
        629 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
        630 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
        631 => x"29292929",		-- colors: 41, 41, 41, 41
        632 => x"29292929",		-- colors: 41, 41, 41, 41
        633 => x"2A292929",		-- colors: 42, 41, 41, 41
        634 => x"2929292A",		-- colors: 41, 41, 41, 42
        635 => x"29292929",		-- colors: 41, 41, 41, 41
        636 => x"29292929",		-- colors: 41, 41, 41, 41
        637 => x"2A292929",		-- colors: 42, 41, 41, 41
        638 => x"2929292A",		-- colors: 41, 41, 41, 42

                --  sprite 6
        639 => x"29292929",		-- colors: 41, 41, 41, 41
        640 => x"29292929",		-- colors: 41, 41, 41, 41
        641 => x"29292929",		-- colors: 41, 41, 41, 41
        642 => x"29292929",		-- colors: 41, 41, 41, 41
        643 => x"29292929",		-- colors: 41, 41, 41, 41
        644 => x"29292929",		-- colors: 41, 41, 41, 41
        645 => x"29292929",		-- colors: 41, 41, 41, 41
        646 => x"29292929",		-- colors: 41, 41, 41, 41
        647 => x"29292929",		-- colors: 41, 41, 41, 41
        648 => x"29292929",		-- colors: 41, 41, 41, 41
        649 => x"29292929",		-- colors: 41, 41, 41, 41
        650 => x"29292929",		-- colors: 41, 41, 41, 41
        651 => x"29292929",		-- colors: 41, 41, 41, 41
        652 => x"29292929",		-- colors: 41, 41, 41, 41
        653 => x"29292929",		-- colors: 41, 41, 41, 41
        654 => x"29292929",		-- colors: 41, 41, 41, 41
        655 => x"29292929",		-- colors: 41, 41, 41, 41
        656 => x"29292929",		-- colors: 41, 41, 41, 41
        657 => x"29292929",		-- colors: 41, 41, 41, 41
        658 => x"29292929",		-- colors: 41, 41, 41, 41
        659 => x"29292929",		-- colors: 41, 41, 41, 41
        660 => x"29292929",		-- colors: 41, 41, 41, 41
        661 => x"29292929",		-- colors: 41, 41, 41, 41
        662 => x"29292929",		-- colors: 41, 41, 41, 41
        663 => x"29292929",		-- colors: 41, 41, 41, 41
        664 => x"29292929",		-- colors: 41, 41, 41, 41
        665 => x"29292929",		-- colors: 41, 41, 41, 41
        666 => x"29292929",		-- colors: 41, 41, 41, 41
        667 => x"29292929",		-- colors: 41, 41, 41, 41
        668 => x"29292929",		-- colors: 41, 41, 41, 41
        669 => x"29292929",		-- colors: 41, 41, 41, 41
        670 => x"29292929",		-- colors: 41, 41, 41, 41
        671 => x"29292929",		-- colors: 41, 41, 41, 41
        672 => x"29292929",		-- colors: 41, 41, 41, 41
        673 => x"29292929",		-- colors: 41, 41, 41, 41
        674 => x"29292929",		-- colors: 41, 41, 41, 41
        675 => x"29292929",		-- colors: 41, 41, 41, 41
        676 => x"29292929",		-- colors: 41, 41, 41, 41
        677 => x"29292929",		-- colors: 41, 41, 41, 41
        678 => x"29292929",		-- colors: 41, 41, 41, 41
        679 => x"29292929",		-- colors: 41, 41, 41, 41
        680 => x"29292929",		-- colors: 41, 41, 41, 41
        681 => x"29292929",		-- colors: 41, 41, 41, 41
        682 => x"29292929",		-- colors: 41, 41, 41, 41
        683 => x"29292929",		-- colors: 41, 41, 41, 41
        684 => x"29292929",		-- colors: 41, 41, 41, 41
        685 => x"29292929",		-- colors: 41, 41, 41, 41
        686 => x"29292929",		-- colors: 41, 41, 41, 41
        687 => x"29292929",		-- colors: 41, 41, 41, 41
        688 => x"29292929",		-- colors: 41, 41, 41, 41
        689 => x"29292929",		-- colors: 41, 41, 41, 41
        690 => x"29292929",		-- colors: 41, 41, 41, 41
        691 => x"29292929",		-- colors: 41, 41, 41, 41
        692 => x"29292929",		-- colors: 41, 41, 41, 41
        693 => x"29292929",		-- colors: 41, 41, 41, 41
        694 => x"29292929",		-- colors: 41, 41, 41, 41
        695 => x"29292929",		-- colors: 41, 41, 41, 41
        696 => x"29292929",		-- colors: 41, 41, 41, 41
        697 => x"29292929",		-- colors: 41, 41, 41, 41
        698 => x"29292929",		-- colors: 41, 41, 41, 41
        699 => x"29292929",		-- colors: 41, 41, 41, 41
        700 => x"29292929",		-- colors: 41, 41, 41, 41
        701 => x"29292929",		-- colors: 41, 41, 41, 41
        702 => x"29292929",		-- colors: 41, 41, 41, 41

                --  sprite 7
        703 => x"28282828",		-- colors: 40, 40, 40, 40
        704 => x"28282828",		-- colors: 40, 40, 40, 40
        705 => x"28282828",		-- colors: 40, 40, 40, 40
        706 => x"28282828",		-- colors: 40, 40, 40, 40
        707 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        708 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        709 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        710 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        711 => x"28282929",		-- colors: 40, 40, 41, 41
        712 => x"29292828",		-- colors: 41, 41, 40, 40
        713 => x"28282929",		-- colors: 40, 40, 41, 41
        714 => x"29292828",		-- colors: 41, 41, 40, 40
        715 => x"28292929",		-- colors: 40, 41, 41, 41
        716 => x"29292928",		-- colors: 41, 41, 41, 40
        717 => x"28292929",		-- colors: 40, 41, 41, 41
        718 => x"29292928",		-- colors: 41, 41, 41, 40
        719 => x"28292929",		-- colors: 40, 41, 41, 41
        720 => x"29292928",		-- colors: 41, 41, 41, 40
        721 => x"28292929",		-- colors: 40, 41, 41, 41
        722 => x"29292928",		-- colors: 41, 41, 41, 40
        723 => x"28282929",		-- colors: 40, 40, 41, 41
        724 => x"29292828",		-- colors: 41, 41, 40, 40
        725 => x"28282929",		-- colors: 40, 40, 41, 41
        726 => x"29292828",		-- colors: 41, 41, 40, 40
        727 => x"28282828",		-- colors: 40, 40, 40, 40
        728 => x"28282828",		-- colors: 40, 40, 40, 40
        729 => x"28282828",		-- colors: 40, 40, 40, 40
        730 => x"28282828",		-- colors: 40, 40, 40, 40
        731 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        732 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        733 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        734 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        735 => x"29292929",		-- colors: 41, 41, 41, 41
        736 => x"29292929",		-- colors: 41, 41, 41, 41
        737 => x"2A292929",		-- colors: 42, 41, 41, 41
        738 => x"2929292A",		-- colors: 41, 41, 41, 42
        739 => x"29292929",		-- colors: 41, 41, 41, 41
        740 => x"29292929",		-- colors: 41, 41, 41, 41
        741 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
        742 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
        743 => x"29292929",		-- colors: 41, 41, 41, 41
        744 => x"29292929",		-- colors: 41, 41, 41, 41
        745 => x"2A292929",		-- colors: 42, 41, 41, 41
        746 => x"2929292A",		-- colors: 41, 41, 41, 42
        747 => x"29292929",		-- colors: 41, 41, 41, 41
        748 => x"29292929",		-- colors: 41, 41, 41, 41
        749 => x"2A292929",		-- colors: 42, 41, 41, 41
        750 => x"2929292A",		-- colors: 41, 41, 41, 42
        751 => x"29292929",		-- colors: 41, 41, 41, 41
        752 => x"29292929",		-- colors: 41, 41, 41, 41
        753 => x"2A292929",		-- colors: 42, 41, 41, 41
        754 => x"2929292A",		-- colors: 41, 41, 41, 42
        755 => x"29292929",		-- colors: 41, 41, 41, 41
        756 => x"29292929",		-- colors: 41, 41, 41, 41
        757 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
        758 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
        759 => x"29292929",		-- colors: 41, 41, 41, 41
        760 => x"29292929",		-- colors: 41, 41, 41, 41
        761 => x"2A292929",		-- colors: 42, 41, 41, 41
        762 => x"2929292A",		-- colors: 41, 41, 41, 42
        763 => x"29292929",		-- colors: 41, 41, 41, 41
        764 => x"29292929",		-- colors: 41, 41, 41, 41
        765 => x"2A292929",		-- colors: 42, 41, 41, 41
        766 => x"2929292A",		-- colors: 41, 41, 41, 42

                --  sprite 8
        767 => x"28282828",		-- colors: 40, 40, 40, 40
        768 => x"28282828",		-- colors: 40, 40, 40, 40
        769 => x"28282828",		-- colors: 40, 40, 40, 40
        770 => x"28282828",		-- colors: 40, 40, 40, 40
        771 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        772 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        773 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        774 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        775 => x"28282929",		-- colors: 40, 40, 41, 41
        776 => x"29292828",		-- colors: 41, 41, 40, 40
        777 => x"28282929",		-- colors: 40, 40, 41, 41
        778 => x"29292828",		-- colors: 41, 41, 40, 40
        779 => x"28292929",		-- colors: 40, 41, 41, 41
        780 => x"29292928",		-- colors: 41, 41, 41, 40
        781 => x"28292929",		-- colors: 40, 41, 41, 41
        782 => x"29292928",		-- colors: 41, 41, 41, 40
        783 => x"28292929",		-- colors: 40, 41, 41, 41
        784 => x"29292928",		-- colors: 41, 41, 41, 40
        785 => x"28292929",		-- colors: 40, 41, 41, 41
        786 => x"29292928",		-- colors: 41, 41, 41, 40
        787 => x"28282929",		-- colors: 40, 40, 41, 41
        788 => x"29292828",		-- colors: 41, 41, 40, 40
        789 => x"28282929",		-- colors: 40, 40, 41, 41
        790 => x"29292828",		-- colors: 41, 41, 40, 40
        791 => x"28282828",		-- colors: 40, 40, 40, 40
        792 => x"28282828",		-- colors: 40, 40, 40, 40
        793 => x"28282828",		-- colors: 40, 40, 40, 40
        794 => x"28282828",		-- colors: 40, 40, 40, 40
        795 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        796 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        797 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        798 => x"2B2B2B2B",		-- colors: 43, 43, 43, 43
        799 => x"2A292929",		-- colors: 42, 41, 41, 41
        800 => x"2929292A",		-- colors: 41, 41, 41, 42
        801 => x"29292929",		-- colors: 41, 41, 41, 41
        802 => x"29292929",		-- colors: 41, 41, 41, 41
        803 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
        804 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
        805 => x"29292929",		-- colors: 41, 41, 41, 41
        806 => x"29292929",		-- colors: 41, 41, 41, 41
        807 => x"2A292929",		-- colors: 42, 41, 41, 41
        808 => x"2929292A",		-- colors: 41, 41, 41, 42
        809 => x"29292929",		-- colors: 41, 41, 41, 41
        810 => x"29292929",		-- colors: 41, 41, 41, 41
        811 => x"2A292929",		-- colors: 42, 41, 41, 41
        812 => x"2929292A",		-- colors: 41, 41, 41, 42
        813 => x"29292929",		-- colors: 41, 41, 41, 41
        814 => x"29292929",		-- colors: 41, 41, 41, 41
        815 => x"2A292929",		-- colors: 42, 41, 41, 41
        816 => x"2929292A",		-- colors: 41, 41, 41, 42
        817 => x"29292929",		-- colors: 41, 41, 41, 41
        818 => x"29292929",		-- colors: 41, 41, 41, 41
        819 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
        820 => x"2A2A2A2A",		-- colors: 42, 42, 42, 42
        821 => x"29292929",		-- colors: 41, 41, 41, 41
        822 => x"29292929",		-- colors: 41, 41, 41, 41
        823 => x"2A292929",		-- colors: 42, 41, 41, 41
        824 => x"2929292A",		-- colors: 41, 41, 41, 42
        825 => x"29292929",		-- colors: 41, 41, 41, 41
        826 => x"29292929",		-- colors: 41, 41, 41, 41
        827 => x"2A292929",		-- colors: 42, 41, 41, 41
        828 => x"2929292A",		-- colors: 41, 41, 41, 42
        829 => x"29292929",		-- colors: 41, 41, 41, 41
        830 => x"29292929",		-- colors: 41, 41, 41, 41
				----------------------------------------------------

				--**VATRICE**--


                --  sprite 0
    831 => x"00000000",		-- colors: 35, 35, 35, 35
        832 => x"00000000",		-- colors: 35, 35, 35, 35
        833 => x"00000000",		-- colors: 35, 35, 35, 35
        834 => x"00000000",		-- colors: 35, 35, 35, 35
        835 => x"00000000",		-- colors: 35, 35, 35, 35
        836 => x"00000000",		-- colors: 35, 35, 35, 35
        837 => x"00000000",		-- colors: 35, 35, 35, 35
        838 => x"00000000",		-- colors: 35, 35, 35, 35
        839 => x"00000000",		-- colors: 35, 35, 35, 35
        840 => x"00000000",		-- colors: 35, 35, 35, 35
        841 => x"00000000",		-- colors: 35, 35, 35, 35
        842 => x"00000000",		-- colors: 35, 35, 35, 35
        843 => x"00000000",		-- colors: 35, 35, 35, 35
        844 => x"00000000",		-- colors: 35, 35, 35, 35
        845 => x"00000000",		-- colors: 35, 35, 35, 35
        846 => x"00000000",		-- colors: 35, 35, 35, 35
        847 => x"00000024",		-- colors: 35, 35, 35, 36
        848 => x"24242424",		-- colors: 36, 36, 36, 36
        849 => x"00000000",		-- colors: 35, 35, 35, 35
        850 => x"00000000",		-- colors: 35, 35, 35, 35
        851 => x"00002424",		-- colors: 35, 35, 36, 36
        852 => x"25252525",		-- colors: 37, 37, 37, 37
        853 => x"24240000",		-- colors: 36, 36, 35, 35
        854 => x"00000000",		-- colors: 35, 35, 35, 35
        855 => x"00242425",		-- colors: 35, 36, 36, 37
        856 => x"25252525",		-- colors: 37, 37, 37, 37
        857 => x"25242400",		-- colors: 37, 36, 36, 35
        858 => x"00000000",		-- colors: 35, 35, 35, 35
        859 => x"00242526",		-- colors: 35, 36, 37, 38
        860 => x"24262426",		-- colors: 36, 38, 36, 38
        861 => x"25252424",		-- colors: 37, 37, 36, 36
        862 => x"00240000",		-- colors: 35, 36, 35, 35
        863 => x"00242526",		-- colors: 35, 36, 37, 38
        864 => x"24262426",		-- colors: 36, 38, 36, 38
        865 => x"26252524",		-- colors: 38, 37, 37, 36
        866 => x"00002400",		-- colors: 35, 35, 36, 35
        867 => x"00002425",		-- colors: 35, 35, 36, 37
        868 => x"26262626",		-- colors: 38, 38, 38, 38
        869 => x"26252524",		-- colors: 38, 37, 37, 36
        870 => x"00242400",		-- colors: 35, 36, 36, 35
        871 => x"00242425",		-- colors: 35, 36, 36, 37
        872 => x"26262626",		-- colors: 38, 38, 38, 38
        873 => x"26252524",		-- colors: 38, 37, 37, 36
        874 => x"24242424",		-- colors: 36, 36, 36, 36
        875 => x"24242525",		-- colors: 36, 36, 37, 37
        876 => x"25262626",		-- colors: 37, 38, 38, 38
        877 => x"25252524",		-- colors: 37, 37, 37, 36
        878 => x"24252400",		-- colors: 36, 37, 36, 35
        879 => x"24242525",		-- colors: 36, 36, 37, 37
        880 => x"25252525",		-- colors: 37, 37, 37, 37
        881 => x"25252525",		-- colors: 37, 37, 37, 37
        882 => x"25240000",		-- colors: 37, 36, 35, 35
        883 => x"24242425",		-- colors: 36, 36, 36, 37
        884 => x"25252525",		-- colors: 37, 37, 37, 37
        885 => x"25252524",		-- colors: 37, 37, 37, 36
        886 => x"24000000",		-- colors: 36, 35, 35, 35
        887 => x"00242424",		-- colors: 35, 36, 36, 36
        888 => x"25252525",		-- colors: 37, 37, 37, 37
        889 => x"25242424",		-- colors: 37, 36, 36, 36
        890 => x"00000000",		-- colors: 35, 35, 35, 35
        891 => x"00000024",		-- colors: 35, 35, 35, 36
        892 => x"24242424",		-- colors: 36, 36, 36, 36
        893 => x"24240000",		-- colors: 36, 36, 35, 35
        894 => x"00000000",		-- colors: 35, 35, 35, 35

                --  sprite 1
       895 => x"00000000",		-- colors: 35, 35, 35, 35
        896 => x"00000000",		-- colors: 35, 35, 35, 35
        897 => x"00000000",		-- colors: 35, 35, 35, 35
        898 => x"00000000",		-- colors: 35, 35, 35, 35
        899 => x"00000000",		-- colors: 35, 35, 35, 35
        900 => x"00000000",		-- colors: 35, 35, 35, 35
        901 => x"00000000",		-- colors: 35, 35, 35, 35
        902 => x"00000000",		-- colors: 35, 35, 35, 35
        903 => x"00000000",		-- colors: 35, 35, 35, 35
        904 => x"00000000",		-- colors: 35, 35, 35, 35
        905 => x"00000000",		-- colors: 35, 35, 35, 35
        906 => x"00000000",		-- colors: 35, 35, 35, 35
        907 => x"00000000",		-- colors: 35, 35, 35, 35
        908 => x"00000000",		-- colors: 35, 35, 35, 35
        909 => x"00000000",		-- colors: 35, 35, 35, 35
        910 => x"00000000",		-- colors: 35, 35, 35, 35
        911 => x"00000000",		-- colors: 35, 35, 35, 35
        912 => x"00000000",		-- colors: 35, 35, 35, 35
        913 => x"24242424",		-- colors: 36, 36, 36, 36
        914 => x"24000000",		-- colors: 36, 35, 35, 35
        915 => x"00000000",		-- colors: 35, 35, 35, 35
        916 => x"00002424",		-- colors: 35, 35, 36, 36
        917 => x"25252525",		-- colors: 37, 37, 37, 37
        918 => x"24240000",		-- colors: 36, 36, 35, 35
        919 => x"00000000",		-- colors: 35, 35, 35, 35
        920 => x"00242425",		-- colors: 35, 36, 36, 37
        921 => x"25252525",		-- colors: 37, 37, 37, 37
        922 => x"25242400",		-- colors: 37, 36, 36, 35
        923 => x"00002400",		-- colors: 35, 35, 36, 35
        924 => x"24242525",		-- colors: 36, 36, 37, 37
        925 => x"26242624",		-- colors: 38, 36, 38, 36
        926 => x"26252400",		-- colors: 38, 37, 36, 35
        927 => x"00240000",		-- colors: 35, 36, 35, 35
        928 => x"24252526",		-- colors: 36, 37, 37, 38
        929 => x"26242624",		-- colors: 38, 36, 38, 36
        930 => x"26252400",		-- colors: 38, 37, 36, 35
        931 => x"00242400",		-- colors: 35, 36, 36, 35
        932 => x"24252526",		-- colors: 36, 37, 37, 38
        933 => x"26262626",		-- colors: 38, 38, 38, 38
        934 => x"25240000",		-- colors: 37, 36, 35, 35
        935 => x"24242424",		-- colors: 36, 36, 36, 36
        936 => x"24252526",		-- colors: 36, 37, 37, 38
        937 => x"26262626",		-- colors: 38, 38, 38, 38
        938 => x"25242400",		-- colors: 37, 36, 36, 35
        939 => x"00242524",		-- colors: 35, 36, 37, 36
        940 => x"24252525",		-- colors: 36, 37, 37, 37
        941 => x"26262625",		-- colors: 38, 38, 38, 37
        942 => x"25252424",		-- colors: 37, 37, 36, 36
        943 => x"00002425",		-- colors: 35, 35, 36, 37
        944 => x"25252525",		-- colors: 37, 37, 37, 37
        945 => x"25252525",		-- colors: 37, 37, 37, 37
        946 => x"25252424",		-- colors: 37, 37, 36, 36
        947 => x"00000024",		-- colors: 35, 35, 35, 36
        948 => x"24252525",		-- colors: 36, 37, 37, 37
        949 => x"25252525",		-- colors: 37, 37, 37, 37
        950 => x"25242424",		-- colors: 37, 36, 36, 36
        951 => x"00000000",		-- colors: 35, 35, 35, 35
        952 => x"24242425",		-- colors: 36, 36, 36, 37
        953 => x"25252525",		-- colors: 37, 37, 37, 37
        954 => x"24242400",		-- colors: 36, 36, 36, 35
        955 => x"00000000",		-- colors: 35, 35, 35, 35
        956 => x"00002424",		-- colors: 35, 35, 36, 36
        957 => x"24242424",		-- colors: 36, 36, 36, 36
        958 => x"24000000",		-- colors: 36, 35, 35, 35

				--**majmun1**--

                --  sprite 0
        959 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        960 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        961 => x"2C2C2D2D",		-- colors: 44, 44, 45, 45
        962 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        963 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        964 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        965 => x"2C2C2C2D",		-- colors: 44, 44, 44, 45
        966 => x"2D2D2E2D",		-- colors: 45, 45, 46, 45
        967 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        968 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        969 => x"2C2C2C2D",		-- colors: 44, 44, 44, 45
        970 => x"2D2D2D2E",		-- colors: 45, 45, 45, 46
        971 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        972 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        973 => x"2C2C2C2D",		-- colors: 44, 44, 44, 45
        974 => x"2D2D2D2E",		-- colors: 45, 45, 45, 46
        975 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        976 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        977 => x"2C2C2C2E",		-- colors: 44, 44, 44, 46
        978 => x"2D2D2E2D",		-- colors: 45, 45, 46, 45
        979 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        980 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        981 => x"2C2C2E2D",		-- colors: 44, 44, 46, 45
        982 => x"2D2D2D2E",		-- colors: 45, 45, 45, 46
        983 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        984 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        985 => x"2C2E2D2D",		-- colors: 44, 46, 45, 45
        986 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        987 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        988 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        989 => x"2E2D2D2D",		-- colors: 46, 45, 45, 45
        990 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        991 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        992 => x"2C2C2C2E",		-- colors: 44, 44, 44, 46
        993 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        994 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        995 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        996 => x"2C2C2C2E",		-- colors: 44, 44, 44, 46
        997 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        998 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        999 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1000 => x"2C2C2C2E",		-- colors: 44, 44, 44, 46
        1001 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1002 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1003 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1004 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1005 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1006 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1007 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1008 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1009 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1010 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1011 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1012 => x"2C2C2E2D",		-- colors: 44, 44, 46, 45
        1013 => x"2E2E2D2D",		-- colors: 46, 46, 45, 45
        1014 => x"2D2E2E2D",		-- colors: 45, 46, 46, 45
        1015 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1016 => x"2C2E2D2E",		-- colors: 44, 46, 45, 46
        1017 => x"2E2D2E2E",		-- colors: 46, 45, 46, 46
        1018 => x"2E2E2D2E",		-- colors: 46, 46, 45, 46
        1019 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1020 => x"2E2D2E2E",		-- colors: 46, 45, 46, 46
        1021 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        1022 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46

                --  sprite 1
        1023 => x"2D2E2D2E",		-- colors: 45, 46, 45, 46
        1024 => x"2D2E2D2D",		-- colors: 45, 46, 45, 45
        1025 => x"2D2D2E2E",		-- colors: 45, 45, 46, 46
        1026 => x"2E2E2E2D",		-- colors: 46, 46, 46, 45
        1027 => x"2D2D2E2E",		-- colors: 45, 45, 46, 46
        1028 => x"2E2E2E2D",		-- colors: 46, 46, 46, 45
        1029 => x"2D2E2E2E",		-- colors: 45, 46, 46, 46
        1030 => x"2D2E2D2D",		-- colors: 45, 46, 45, 45
        1031 => x"2D2E2E2E",		-- colors: 45, 46, 46, 46
        1032 => x"2E2E2E2D",		-- colors: 46, 46, 46, 45
        1033 => x"2D2E2E2E",		-- colors: 45, 46, 46, 46
        1034 => x"2E2D2D2D",		-- colors: 46, 45, 45, 45
        1035 => x"2D2E2E2D",		-- colors: 45, 46, 46, 45
        1036 => x"2E2E2E2D",		-- colors: 46, 46, 46, 45
        1037 => x"2D2E2E2E",		-- colors: 45, 46, 46, 46
        1038 => x"2D2E2D2D",		-- colors: 45, 46, 45, 45
        1039 => x"2D2E2E2E",		-- colors: 45, 46, 46, 46
        1040 => x"2E2E2D2E",		-- colors: 46, 46, 45, 46
        1041 => x"2E2D2E2E",		-- colors: 46, 45, 46, 46
        1042 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        1043 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1044 => x"2D2D2E2E",		-- colors: 45, 45, 46, 46
        1045 => x"2E2E2D2E",		-- colors: 46, 46, 45, 46
        1046 => x"2E2E2E2D",		-- colors: 46, 46, 46, 45
        1047 => x"2D2D2D2E",		-- colors: 45, 45, 45, 46
        1048 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        1049 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        1050 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1051 => x"2D2D2E2E",		-- colors: 45, 45, 46, 46
        1052 => x"2D2D2D2E",		-- colors: 45, 45, 45, 46
        1053 => x"2D2D2E2D",		-- colors: 45, 45, 46, 45
        1054 => x"2E2E2D2D",		-- colors: 46, 46, 45, 45
        1055 => x"2D2D2D2E",		-- colors: 45, 45, 45, 46
        1056 => x"2E2D2E2D",		-- colors: 46, 45, 46, 45
        1057 => x"2E2D2D2E",		-- colors: 46, 45, 45, 46
        1058 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1059 => x"2D2D2E2D",		-- colors: 45, 45, 46, 45
        1060 => x"2D2E2D2E",		-- colors: 45, 46, 45, 46
        1061 => x"2D2D2E2D",		-- colors: 45, 45, 46, 45
        1062 => x"2D2E2D2D",		-- colors: 45, 46, 45, 45
        1063 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1064 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1065 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1066 => x"2C2C2D2D",		-- colors: 44, 44, 45, 45
        1067 => x"2D2D2D2C",		-- colors: 45, 45, 45, 44
        1068 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1069 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1070 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1071 => x"2D2D2C2C",		-- colors: 45, 45, 44, 44
        1072 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1073 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1074 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1075 => x"2E2C2C2C",		-- colors: 46, 44, 44, 44
        1076 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1077 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1078 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1079 => x"2E2C2C2C",		-- colors: 46, 44, 44, 44
        1080 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1081 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1082 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1083 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1084 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1085 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1086 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44

                --  sprite 2
        1087 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1088 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1089 => x"2D2D2C2C",		-- colors: 45, 45, 44, 44
        1090 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1091 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1092 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1093 => x"2D2C2C2C",		-- colors: 45, 44, 44, 44
        1094 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1095 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1096 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1097 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1098 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1099 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1100 => x"2D2C2C2C",		-- colors: 45, 44, 44, 44
        1101 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1102 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1103 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1104 => x"2D2E2E2C",		-- colors: 45, 46, 46, 44
        1105 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1106 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1107 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1108 => x"2D2D2D2E",		-- colors: 45, 45, 45, 46
        1109 => x"2E2C2C2C",		-- colors: 46, 44, 44, 44
        1110 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1111 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1112 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1113 => x"2D2E2C2C",		-- colors: 45, 46, 44, 44
        1114 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1115 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1116 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1117 => x"2D2E2C2C",		-- colors: 45, 46, 44, 44
        1118 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1119 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1120 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1121 => x"2D2E2C2C",		-- colors: 45, 46, 44, 44
        1122 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1123 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1124 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1125 => x"2D2E2C2C",		-- colors: 45, 46, 44, 44
        1126 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1127 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1128 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1129 => x"2D2D2D2C",		-- colors: 45, 45, 45, 44
        1130 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1131 => x"2C2C2D2D",		-- colors: 44, 44, 45, 45
        1132 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1133 => x"2D2D2E2E",		-- colors: 45, 45, 46, 46
        1134 => x"2E2C2C2C",		-- colors: 46, 44, 44, 44
        1135 => x"2C2C2C2D",		-- colors: 44, 44, 44, 45
        1136 => x"2D2D2D2E",		-- colors: 45, 45, 45, 46
        1137 => x"2E2E2D2E",		-- colors: 46, 46, 45, 46
        1138 => x"2E2E2C2C",		-- colors: 46, 46, 44, 44
        1139 => x"2C2C2C2E",		-- colors: 44, 44, 44, 46
        1140 => x"2E2E2E2D",		-- colors: 46, 46, 46, 45
        1141 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        1142 => x"2E2E2C2C",		-- colors: 46, 46, 44, 44
        1143 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1144 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1145 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1146 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1147 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1148 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1149 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1150 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44

                --  sprite 3
        1151 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1152 => x"2C2C0000",		-- colors: 44, 44, 46, 46
        1153 => x"00002C2C",		-- colors: 46, 46, 44, 44
        1154 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1155 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1156 => x"00000000",		-- colors: 46, 46, 46, 46
        1157 => x"2D2E2E2C",		-- colors: 45, 46, 46, 44
        1158 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1159 => x"2C2C2E2E",		-- colors: 44, 44, 46, 46
        1160 => x"00000000",		-- colors: 46, 45, 46, 46
        1161 => x"2E2D2E2E",		-- colors: 46, 45, 46, 46
        1162 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1163 => x"2C2C2E2E",		-- colors: 44, 44, 46, 46
        1164 => x"00000000",		-- colors: 46, 46, 45, 46
        1165 => x"2D2D2D2C",		-- colors: 45, 45, 45, 44
        1166 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1167 => x"2C2D2E2D",		-- colors: 44, 45, 46, 45
        1168 => x"00000000",		-- colors: 46, 46, 46, 45
        1169 => x"2E2E2E2C",		-- colors: 46, 46, 46, 44
        1170 => x"2C2C2C2E",		-- colors: 44, 44, 44, 46
        1171 => x"2C2D2D2D",		-- colors: 44, 45, 45, 45
        1172 => x"2D2E2E2E",		-- colors: 45, 46, 46, 46
        1173 => x"2E2E2C2C",		-- colors: 46, 46, 44, 44
        1174 => x"2C2C2E2E",		-- colors: 44, 44, 46, 46
        1175 => x"2C2D2D2D",		-- colors: 44, 45, 45, 45
        1176 => x"2D2D2D2C",		-- colors: 45, 45, 45, 44
        1177 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1178 => x"2C2D2E2E",		-- colors: 44, 45, 46, 46
        1179 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1180 => x"2D2D2E2D",		-- colors: 45, 45, 46, 45
        1181 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1182 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1183 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1184 => x"2D2E2D2D",		-- colors: 45, 46, 45, 45
        1185 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1186 => x"2D2D2D2E",		-- colors: 45, 45, 45, 46
        1187 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1188 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1189 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1190 => x"2D2D2D2E",		-- colors: 45, 45, 45, 46
        1191 => x"2C2D2D2D",		-- colors: 44, 45, 45, 45
        1192 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1193 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1194 => x"2D2D2D2E",		-- colors: 45, 45, 45, 46
        1195 => x"2C2C2D2D",		-- colors: 44, 44, 45, 45
        1196 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1197 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1198 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1199 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1200 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1201 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1202 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1203 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1204 => x"2C2D2D2D",		-- colors: 44, 45, 45, 45
        1205 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1206 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1207 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1208 => x"2C2C2C2D",		-- colors: 44, 44, 44, 45
        1209 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1210 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1211 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1212 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1213 => x"2C2D2D2D",		-- colors: 44, 45, 45, 45
        1214 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45

                --  sprite 4
        1215 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1216 => x"2C2D2D2D",		-- colors: 44, 45, 45, 45
        1217 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1218 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1219 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1220 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1221 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1222 => x"2D2C2C2C",		-- colors: 45, 44, 44, 44
        1223 => x"2C2C2C2D",		-- colors: 44, 44, 44, 45
        1224 => x"2D2E2E2D",		-- colors: 45, 46, 46, 45
        1225 => x"2D2D2E2E",		-- colors: 45, 45, 46, 46
        1226 => x"2D2D2C2C",		-- colors: 45, 45, 44, 44
        1227 => x"2C2C2D2D",		-- colors: 44, 44, 45, 45
        1228 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        1229 => x"2D2E2E2E",		-- colors: 45, 46, 46, 46
        1230 => x"2E2D2D2C",		-- colors: 46, 45, 45, 44
        1231 => x"2E2D2D2E",		-- colors: 46, 45, 45, 46
        1232 => x"2E2E2F2F",		-- colors: 46, 46, 47, 47
        1233 => x"2E2F2F2E",		-- colors: 46, 47, 47, 46
        1234 => x"2E2E2D2E",		-- colors: 46, 46, 45, 46
        1235 => x"2E2D2D2D",		-- colors: 46, 45, 45, 45
        1236 => x"2E2E2F2C",		-- colors: 46, 46, 47, 44
        1237 => x"2E2C2F2E",		-- colors: 46, 44, 47, 46
        1238 => x"2E2D2D2E",		-- colors: 46, 45, 45, 46
        1239 => x"2E2D2D2D",		-- colors: 46, 45, 45, 45
        1240 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        1241 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        1242 => x"2E2D2D2E",		-- colors: 46, 45, 45, 46
        1243 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        1244 => x"2E2E2E2D",		-- colors: 46, 46, 46, 45
        1245 => x"2D2D2E2E",		-- colors: 45, 45, 46, 46
        1246 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        1247 => x"2E2E2F2F",		-- colors: 46, 46, 47, 47
        1248 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        1249 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        1250 => x"2E2F2F2E",		-- colors: 46, 47, 47, 46
        1251 => x"2E2F2F2F",		-- colors: 46, 47, 47, 47
        1252 => x"2D2F2F2F",		-- colors: 45, 47, 47, 47
        1253 => x"2D2F2F2F",		-- colors: 45, 47, 47, 47
        1254 => x"2D2F2F2F",		-- colors: 45, 47, 47, 47
        1255 => x"2E2D2F2D",		-- colors: 46, 45, 47, 45
        1256 => x"2D2D2F2D",		-- colors: 45, 45, 47, 45
        1257 => x"2D2D2F2D",		-- colors: 45, 45, 47, 45
        1258 => x"2D2D2F2D",		-- colors: 45, 45, 47, 45
        1259 => x"2E2E2F2F",		-- colors: 46, 46, 47, 47
        1260 => x"2D2F2F2F",		-- colors: 45, 47, 47, 47
        1261 => x"2D2F2F2F",		-- colors: 45, 47, 47, 47
        1262 => x"2D2F2F2E",		-- colors: 45, 47, 47, 46
        1263 => x"2D2E2E2E",		-- colors: 45, 46, 46, 46
        1264 => x"2E2F2F2F",		-- colors: 46, 47, 47, 47
        1265 => x"2F2F2F2F",		-- colors: 47, 47, 47, 47
        1266 => x"2E2E2E2D",		-- colors: 46, 46, 46, 45
        1267 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1268 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        1269 => x"2E2E2E2E",		-- colors: 46, 46, 46, 46
        1270 => x"2E2D2D2D",		-- colors: 46, 45, 45, 45
        1271 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1272 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1273 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1274 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1275 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1276 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1277 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1278 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45

                --  sprite 5
        1279 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1280 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1281 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1282 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1283 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1284 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1285 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1286 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1287 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1288 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1289 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1290 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1291 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1292 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1293 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1294 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1295 => x"2E2C2C2C",		-- colors: 46, 44, 44, 44
        1296 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1297 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1298 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1299 => x"2E2E2C2C",		-- colors: 46, 46, 44, 44
        1300 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1301 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1302 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1303 => x"2E2E2C2C",		-- colors: 46, 46, 44, 44
        1304 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1305 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1306 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1307 => x"2D2D2D2E",		-- colors: 45, 45, 45, 46
        1308 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1309 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1310 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1311 => x"2E2D2D2D",		-- colors: 46, 45, 45, 45
        1312 => x"2E2E2C2C",		-- colors: 46, 46, 44, 44
        1313 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1314 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1315 => x"2E2D2D2D",		-- colors: 46, 45, 45, 45
        1316 => x"2D2D2E2C",		-- colors: 45, 45, 46, 44
        1317 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1318 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1319 => x"2E2D2D2D",		-- colors: 46, 45, 45, 45
        1320 => x"2D2D2D2E",		-- colors: 45, 45, 45, 46
        1321 => x"2E2C2C2C",		-- colors: 46, 44, 44, 44
        1322 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1323 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1324 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1325 => x"2D2E2C2C",		-- colors: 45, 46, 44, 44
        1326 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1327 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1328 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1329 => x"2D2D2E2C",		-- colors: 45, 45, 46, 44
        1330 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1331 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1332 => x"2E2D2D2D",		-- colors: 46, 45, 45, 45
        1333 => x"2D2D2D2C",		-- colors: 45, 45, 45, 44
        1334 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1335 => x"2D2D2D2E",		-- colors: 45, 45, 45, 46
        1336 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1337 => x"2D2D2D2C",		-- colors: 45, 45, 45, 44
        1338 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
        1339 => x"2E2E2E2D",		-- colors: 46, 46, 46, 45
        1340 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
        1341 => x"2D2D2D2C",		-- colors: 45, 45, 45, 44
        1342 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44

				--**majmun2**

                --  sprite 0
        1343 => x"30303030",		-- colors: 48, 48, 48, 48
        1344 => x"30303030",		-- colors: 48, 48, 48, 48
        1345 => x"30303030",		-- colors: 48, 48, 48, 48
        1346 => x"30303030",		-- colors: 48, 48, 48, 48
        1347 => x"30303030",		-- colors: 48, 48, 48, 48
        1348 => x"30303030",		-- colors: 48, 48, 48, 48
        1349 => x"30303030",		-- colors: 48, 48, 48, 48
        1350 => x"30303030",		-- colors: 48, 48, 48, 48
        1351 => x"30303030",		-- colors: 48, 48, 48, 48
        1352 => x"30303030",		-- colors: 48, 48, 48, 48
        1353 => x"30303030",		-- colors: 48, 48, 48, 48
        1354 => x"30303030",		-- colors: 48, 48, 48, 48
        1355 => x"30303030",		-- colors: 48, 48, 48, 48
        1356 => x"30303030",		-- colors: 48, 48, 48, 48
        1357 => x"30303030",		-- colors: 48, 48, 48, 48
        1358 => x"30303030",		-- colors: 48, 48, 48, 48
        1359 => x"30303030",		-- colors: 48, 48, 48, 48
        1360 => x"30303030",		-- colors: 48, 48, 48, 48
        1361 => x"30303030",		-- colors: 48, 48, 48, 48
        1362 => x"30303032",		-- colors: 48, 48, 48, 50
        1363 => x"30303030",		-- colors: 48, 48, 48, 48
        1364 => x"30303030",		-- colors: 48, 48, 48, 48
        1365 => x"30303030",		-- colors: 48, 48, 48, 48
        1366 => x"30303232",		-- colors: 48, 48, 50, 50
        1367 => x"30303030",		-- colors: 48, 48, 48, 48
        1368 => x"30303030",		-- colors: 48, 48, 48, 48
        1369 => x"30303030",		-- colors: 48, 48, 48, 48
        1370 => x"30303232",		-- colors: 48, 48, 50, 50
        1371 => x"30303030",		-- colors: 48, 48, 48, 48
        1372 => x"30303030",		-- colors: 48, 48, 48, 48
        1373 => x"30303030",		-- colors: 48, 48, 48, 48
        1374 => x"32313131",		-- colors: 50, 49, 49, 49
        1375 => x"30303030",		-- colors: 48, 48, 48, 48
        1376 => x"30303030",		-- colors: 48, 48, 48, 48
        1377 => x"30303232",		-- colors: 48, 48, 50, 50
        1378 => x"31313132",		-- colors: 49, 49, 49, 50
        1379 => x"30303030",		-- colors: 48, 48, 48, 48
        1380 => x"30303030",		-- colors: 48, 48, 48, 48
        1381 => x"30323131",		-- colors: 48, 50, 49, 49
        1382 => x"31313132",		-- colors: 49, 49, 49, 50
        1383 => x"30303030",		-- colors: 48, 48, 48, 48
        1384 => x"30303032",		-- colors: 48, 48, 48, 50
        1385 => x"32313131",		-- colors: 50, 49, 49, 49
        1386 => x"31313132",		-- colors: 49, 49, 49, 50
        1387 => x"30303030",		-- colors: 48, 48, 48, 48
        1388 => x"30303231",		-- colors: 48, 48, 50, 49
        1389 => x"31313131",		-- colors: 49, 49, 49, 49
        1390 => x"31313131",		-- colors: 49, 49, 49, 49
        1391 => x"30303030",		-- colors: 48, 48, 48, 48
        1392 => x"30323131",		-- colors: 48, 50, 49, 49
        1393 => x"31313131",		-- colors: 49, 49, 49, 49
        1394 => x"31313131",		-- colors: 49, 49, 49, 49
        1395 => x"30303030",		-- colors: 48, 48, 48, 48
        1396 => x"30313131",		-- colors: 48, 49, 49, 49
        1397 => x"31313132",		-- colors: 49, 49, 49, 50
        1398 => x"31313131",		-- colors: 49, 49, 49, 49
        1399 => x"30303030",		-- colors: 48, 48, 48, 48
        1400 => x"30313131",		-- colors: 48, 49, 49, 49
        1401 => x"31313131",		-- colors: 49, 49, 49, 49
        1402 => x"32313131",		-- colors: 50, 49, 49, 49
        1403 => x"30303030",		-- colors: 48, 48, 48, 48
        1404 => x"30313131",		-- colors: 48, 49, 49, 49
        1405 => x"31313131",		-- colors: 49, 49, 49, 49
        1406 => x"31323232",		-- colors: 49, 50, 50, 50

                --  sprite 1
        1407 => x"30303030",		-- colors: 48, 48, 48, 48
        1408 => x"31313131",		-- colors: 49, 49, 49, 49
        1409 => x"31313130",		-- colors: 49, 49, 49, 48
        1410 => x"30303030",		-- colors: 48, 48, 48, 48
        1411 => x"30303031",		-- colors: 48, 48, 48, 49
        1412 => x"31313131",		-- colors: 49, 49, 49, 49
        1413 => x"31313131",		-- colors: 49, 49, 49, 49
        1414 => x"30303030",		-- colors: 48, 48, 48, 48
        1415 => x"30303131",		-- colors: 48, 48, 49, 49
        1416 => x"32323131",		-- colors: 50, 50, 49, 49
        1417 => x"31323231",		-- colors: 49, 50, 50, 49
        1418 => x"31303030",		-- colors: 49, 48, 48, 48
        1419 => x"30313132",		-- colors: 48, 49, 49, 50
        1420 => x"32323231",		-- colors: 50, 50, 50, 49
        1421 => x"32323232",		-- colors: 50, 50, 50, 50
        1422 => x"31313030",		-- colors: 49, 49, 48, 48
        1423 => x"32313232",		-- colors: 50, 49, 50, 50
        1424 => x"32333332",		-- colors: 50, 51, 51, 50
        1425 => x"33333232",		-- colors: 51, 51, 50, 50
        1426 => x"32313132",		-- colors: 50, 49, 49, 50
        1427 => x"32313132",		-- colors: 50, 49, 49, 50
        1428 => x"32333032",		-- colors: 50, 51, 48, 50
        1429 => x"30333232",		-- colors: 48, 51, 50, 50
        1430 => x"31313132",		-- colors: 49, 49, 49, 50
        1431 => x"32313132",		-- colors: 50, 49, 49, 50
        1432 => x"32323232",		-- colors: 50, 50, 50, 50
        1433 => x"32323232",		-- colors: 50, 50, 50, 50
        1434 => x"31313132",		-- colors: 49, 49, 49, 50
        1435 => x"32323232",		-- colors: 50, 50, 50, 50
        1436 => x"32323131",		-- colors: 50, 50, 49, 49
        1437 => x"31323232",		-- colors: 49, 50, 50, 50
        1438 => x"32323232",		-- colors: 50, 50, 50, 50
        1439 => x"32333332",		-- colors: 50, 51, 51, 50
        1440 => x"32323232",		-- colors: 50, 50, 50, 50
        1441 => x"32323232",		-- colors: 50, 50, 50, 50
        1442 => x"33333232",		-- colors: 51, 51, 50, 50
        1443 => x"33333331",		-- colors: 51, 51, 51, 49
        1444 => x"33333331",		-- colors: 51, 51, 51, 49
        1445 => x"33333331",		-- colors: 51, 51, 51, 49
        1446 => x"33333332",		-- colors: 51, 51, 51, 50
        1447 => x"31333131",		-- colors: 49, 51, 49, 49
        1448 => x"31333131",		-- colors: 49, 51, 49, 49
        1449 => x"31333131",		-- colors: 49, 51, 49, 49
        1450 => x"31333132",		-- colors: 49, 51, 49, 50
        1451 => x"32333331",		-- colors: 50, 51, 51, 49
        1452 => x"33333331",		-- colors: 51, 51, 51, 49
        1453 => x"33333331",		-- colors: 51, 51, 51, 49
        1454 => x"33333232",		-- colors: 51, 51, 50, 50
        1455 => x"31323232",		-- colors: 49, 50, 50, 50
        1456 => x"33333333",		-- colors: 51, 51, 51, 51
        1457 => x"33333332",		-- colors: 51, 51, 51, 50
        1458 => x"32323231",		-- colors: 50, 50, 50, 49
        1459 => x"31313132",		-- colors: 49, 49, 49, 50
        1460 => x"32323232",		-- colors: 50, 50, 50, 50
        1461 => x"32323232",		-- colors: 50, 50, 50, 50
        1462 => x"31313131",		-- colors: 49, 49, 49, 49
        1463 => x"31313131",		-- colors: 49, 49, 49, 49
        1464 => x"31313131",		-- colors: 49, 49, 49, 49
        1465 => x"31313131",		-- colors: 49, 49, 49, 49
        1466 => x"31313131",		-- colors: 49, 49, 49, 49
        1467 => x"31313131",		-- colors: 49, 49, 49, 49
        1468 => x"31313131",		-- colors: 49, 49, 49, 49
        1469 => x"31313131",		-- colors: 49, 49, 49, 49
        1470 => x"31313131",		-- colors: 49, 49, 49, 49

                --  sprite 2
        1471 => x"30303030",		-- colors: 48, 48, 48, 48
        1472 => x"30303232",		-- colors: 48, 48, 50, 50
        1473 => x"32323030",		-- colors: 50, 50, 48, 48
        1474 => x"30303030",		-- colors: 48, 48, 48, 48
        1475 => x"30303030",		-- colors: 48, 48, 48, 48
        1476 => x"30323231",		-- colors: 48, 50, 50, 49
        1477 => x"32323232",		-- colors: 50, 50, 50, 50
        1478 => x"30303030",		-- colors: 48, 48, 48, 48
        1479 => x"30303030",		-- colors: 48, 48, 48, 48
        1480 => x"32323132",		-- colors: 50, 50, 49, 50
        1481 => x"32323132",		-- colors: 50, 50, 49, 50
        1482 => x"32323030",		-- colors: 50, 50, 48, 48
        1483 => x"30303030",		-- colors: 48, 48, 48, 48
        1484 => x"30313131",		-- colors: 48, 49, 49, 49
        1485 => x"32313232",		-- colors: 50, 49, 50, 50
        1486 => x"32323030",		-- colors: 50, 50, 48, 48
        1487 => x"32303030",		-- colors: 50, 48, 48, 48
        1488 => x"30323232",		-- colors: 48, 50, 50, 50
        1489 => x"31323232",		-- colors: 49, 50, 50, 50
        1490 => x"31323130",		-- colors: 49, 50, 49, 48
        1491 => x"32323030",		-- colors: 50, 50, 48, 48
        1492 => x"30303232",		-- colors: 48, 48, 50, 50
        1493 => x"32323231",		-- colors: 50, 50, 50, 49
        1494 => x"31313130",		-- colors: 49, 49, 49, 48
        1495 => x"32323130",		-- colors: 50, 50, 49, 48
        1496 => x"30303030",		-- colors: 48, 48, 48, 48
        1497 => x"30313131",		-- colors: 48, 49, 49, 49
        1498 => x"31313130",		-- colors: 49, 49, 49, 48
        1499 => x"31313131",		-- colors: 49, 49, 49, 49
        1500 => x"31313131",		-- colors: 49, 49, 49, 49
        1501 => x"31323131",		-- colors: 49, 50, 49, 49
        1502 => x"31313131",		-- colors: 49, 49, 49, 49
        1503 => x"32313131",		-- colors: 50, 49, 49, 49
        1504 => x"31313131",		-- colors: 49, 49, 49, 49
        1505 => x"31313231",		-- colors: 49, 49, 50, 49
        1506 => x"31313131",		-- colors: 49, 49, 49, 49
        1507 => x"32313131",		-- colors: 50, 49, 49, 49
        1508 => x"31313131",		-- colors: 49, 49, 49, 49
        1509 => x"31313131",		-- colors: 49, 49, 49, 49
        1510 => x"31313131",		-- colors: 49, 49, 49, 49
        1511 => x"32313131",		-- colors: 50, 49, 49, 49
        1512 => x"31313131",		-- colors: 49, 49, 49, 49
        1513 => x"31313131",		-- colors: 49, 49, 49, 49
        1514 => x"31313130",		-- colors: 49, 49, 49, 48
        1515 => x"31313131",		-- colors: 49, 49, 49, 49
        1516 => x"31313131",		-- colors: 49, 49, 49, 49
        1517 => x"31313131",		-- colors: 49, 49, 49, 49
        1518 => x"31313030",		-- colors: 49, 49, 48, 48
        1519 => x"31313131",		-- colors: 49, 49, 49, 49
        1520 => x"31313131",		-- colors: 49, 49, 49, 49
        1521 => x"31313131",		-- colors: 49, 49, 49, 49
        1522 => x"30303030",		-- colors: 48, 48, 48, 48
        1523 => x"31313131",		-- colors: 49, 49, 49, 49
        1524 => x"31313131",		-- colors: 49, 49, 49, 49
        1525 => x"31313130",		-- colors: 49, 49, 49, 48
        1526 => x"30303030",		-- colors: 48, 48, 48, 48
        1527 => x"31313131",		-- colors: 49, 49, 49, 49
        1528 => x"31313131",		-- colors: 49, 49, 49, 49
        1529 => x"31303030",		-- colors: 49, 48, 48, 48
        1530 => x"30303030",		-- colors: 48, 48, 48, 48
        1531 => x"31313131",		-- colors: 49, 49, 49, 49
        1532 => x"31313130",		-- colors: 49, 49, 49, 48
        1533 => x"30303030",		-- colors: 48, 48, 48, 48
        1534 => x"30303030",		-- colors: 48, 48, 48, 48

                --  sprite 3
        1535 => x"30303030",		-- colors: 48, 48, 48, 48
        1536 => x"30303131",		-- colors: 48, 48, 49, 49
        1537 => x"31313131",		-- colors: 49, 49, 49, 49
        1538 => x"31313131",		-- colors: 49, 49, 49, 49
        1539 => x"30303030",		-- colors: 48, 48, 48, 48
        1540 => x"30303031",		-- colors: 48, 48, 48, 49
        1541 => x"31313131",		-- colors: 49, 49, 49, 49
        1542 => x"31313131",		-- colors: 49, 49, 49, 49
        1543 => x"30303030",		-- colors: 48, 48, 48, 48
        1544 => x"30303030",		-- colors: 48, 48, 48, 48
        1545 => x"31313131",		-- colors: 49, 49, 49, 49
        1546 => x"31313131",		-- colors: 49, 49, 49, 49
        1547 => x"30303030",		-- colors: 48, 48, 48, 48
        1548 => x"30303030",		-- colors: 48, 48, 48, 48
        1549 => x"30303031",		-- colors: 48, 48, 48, 49
        1550 => x"31313131",		-- colors: 49, 49, 49, 49
        1551 => x"30303030",		-- colors: 48, 48, 48, 48
        1552 => x"30303030",		-- colors: 48, 48, 48, 48
        1553 => x"30323231",		-- colors: 48, 50, 50, 49
        1554 => x"31313131",		-- colors: 49, 49, 49, 49
        1555 => x"30303030",		-- colors: 48, 48, 48, 48
        1556 => x"30303032",		-- colors: 48, 48, 48, 50
        1557 => x"32313131",		-- colors: 50, 49, 49, 49
        1558 => x"31313131",		-- colors: 49, 49, 49, 49
        1559 => x"30303030",		-- colors: 48, 48, 48, 48
        1560 => x"30303231",		-- colors: 48, 48, 50, 49
        1561 => x"31313131",		-- colors: 49, 49, 49, 49
        1562 => x"31313131",		-- colors: 49, 49, 49, 49
        1563 => x"30303030",		-- colors: 48, 48, 48, 48
        1564 => x"30303231",		-- colors: 48, 48, 50, 49
        1565 => x"31313131",		-- colors: 49, 49, 49, 49
        1566 => x"31313131",		-- colors: 49, 49, 49, 49
        1567 => x"30303030",		-- colors: 48, 48, 48, 48
        1568 => x"30303231",		-- colors: 48, 48, 50, 49
        1569 => x"31313131",		-- colors: 49, 49, 49, 49
        1570 => x"31313131",		-- colors: 49, 49, 49, 49
        1571 => x"30303030",		-- colors: 48, 48, 48, 48
        1572 => x"30303231",		-- colors: 48, 48, 50, 49
        1573 => x"31313131",		-- colors: 49, 49, 49, 49
        1574 => x"31313131",		-- colors: 49, 49, 49, 49
        1575 => x"30303030",		-- colors: 48, 48, 48, 48
        1576 => x"30313131",		-- colors: 48, 49, 49, 49
        1577 => x"31313131",		-- colors: 49, 49, 49, 49
        1578 => x"31313131",		-- colors: 49, 49, 49, 49
        1579 => x"30303032",		-- colors: 48, 48, 48, 50
        1580 => x"32323131",		-- colors: 50, 50, 49, 49
        1581 => x"31313131",		-- colors: 49, 49, 49, 49
        1582 => x"31313030",		-- colors: 49, 49, 48, 48
        1583 => x"30303232",		-- colors: 48, 48, 50, 50
        1584 => x"32313232",		-- colors: 50, 49, 50, 50
        1585 => x"32313131",		-- colors: 50, 49, 49, 49
        1586 => x"31303030",		-- colors: 49, 48, 48, 48
        1587 => x"30303232",		-- colors: 48, 48, 50, 50
        1588 => x"32323232",		-- colors: 50, 50, 50, 50
        1589 => x"31323232",		-- colors: 49, 50, 50, 50
        1590 => x"32303030",		-- colors: 50, 48, 48, 48
        1591 => x"30303030",		-- colors: 48, 48, 48, 48
        1592 => x"30303030",		-- colors: 48, 48, 48, 48
        1593 => x"30303030",		-- colors: 48, 48, 48, 48
        1594 => x"30303030",		-- colors: 48, 48, 48, 48
        1595 => x"30303030",		-- colors: 48, 48, 48, 48
        1596 => x"30303030",		-- colors: 48, 48, 48, 48
        1597 => x"30303030",		-- colors: 48, 48, 48, 48
        1598 => x"30303030",		-- colors: 48, 48, 48, 48

                --  sprite 4
        1599 => x"31323232",		-- colors: 49, 50, 50, 50
        1600 => x"32323131",		-- colors: 50, 50, 49, 49
        1601 => x"31313231",		-- colors: 49, 49, 50, 49
        1602 => x"32313231",		-- colors: 50, 49, 50, 49
        1603 => x"31313231",		-- colors: 49, 49, 50, 49
        1604 => x"32323231",		-- colors: 50, 50, 50, 49
        1605 => x"31323232",		-- colors: 49, 50, 50, 50
        1606 => x"32323131",		-- colors: 50, 50, 49, 49
        1607 => x"31313132",		-- colors: 49, 49, 49, 50
        1608 => x"32323231",		-- colors: 50, 50, 50, 49
        1609 => x"31323232",		-- colors: 49, 50, 50, 50
        1610 => x"32323231",		-- colors: 50, 50, 50, 49
        1611 => x"31313231",		-- colors: 49, 49, 50, 49
        1612 => x"32323231",		-- colors: 50, 50, 50, 49
        1613 => x"31323232",		-- colors: 49, 50, 50, 50
        1614 => x"31323231",		-- colors: 49, 50, 50, 49
        1615 => x"32323232",		-- colors: 50, 50, 50, 50
        1616 => x"32323132",		-- colors: 50, 50, 49, 50
        1617 => x"32313232",		-- colors: 50, 49, 50, 50
        1618 => x"32323231",		-- colors: 50, 50, 50, 49
        1619 => x"31323232",		-- colors: 49, 50, 50, 50
        1620 => x"32313232",		-- colors: 50, 49, 50, 50
        1621 => x"32323131",		-- colors: 50, 50, 49, 49
        1622 => x"31313131",		-- colors: 49, 49, 49, 49
        1623 => x"31313131",		-- colors: 49, 49, 49, 49
        1624 => x"32323232",		-- colors: 50, 50, 50, 50
        1625 => x"32323232",		-- colors: 50, 50, 50, 50
        1626 => x"32313131",		-- colors: 50, 49, 49, 49
        1627 => x"31313232",		-- colors: 49, 49, 50, 50
        1628 => x"31323131",		-- colors: 49, 50, 49, 49
        1629 => x"32313131",		-- colors: 50, 49, 49, 49
        1630 => x"32323131",		-- colors: 50, 50, 49, 49
        1631 => x"31313131",		-- colors: 49, 49, 49, 49
        1632 => x"32313132",		-- colors: 50, 49, 49, 50
        1633 => x"31323132",		-- colors: 49, 50, 49, 50
        1634 => x"32313131",		-- colors: 50, 49, 49, 49
        1635 => x"31313231",		-- colors: 49, 49, 50, 49
        1636 => x"31323131",		-- colors: 49, 50, 49, 49
        1637 => x"32313231",		-- colors: 50, 49, 50, 49
        1638 => x"31323131",		-- colors: 49, 50, 49, 49
        1639 => x"31313030",		-- colors: 49, 49, 48, 48
        1640 => x"30303030",		-- colors: 48, 48, 48, 48
        1641 => x"30303030",		-- colors: 48, 48, 48, 48
        1642 => x"31313131",		-- colors: 49, 49, 49, 49
        1643 => x"30303030",		-- colors: 48, 48, 48, 48
        1644 => x"30303030",		-- colors: 48, 48, 48, 48
        1645 => x"30303030",		-- colors: 48, 48, 48, 48
        1646 => x"30313131",		-- colors: 48, 49, 49, 49
        1647 => x"30303030",		-- colors: 48, 48, 48, 48
        1648 => x"30303030",		-- colors: 48, 48, 48, 48
        1649 => x"30303030",		-- colors: 48, 48, 48, 48
        1650 => x"30303131",		-- colors: 48, 48, 49, 49
        1651 => x"30303030",		-- colors: 48, 48, 48, 48
        1652 => x"30303030",		-- colors: 48, 48, 48, 48
        1653 => x"30303030",		-- colors: 48, 48, 48, 48
        1654 => x"30303032",		-- colors: 48, 48, 48, 50
        1655 => x"30303030",		-- colors: 48, 48, 48, 48
        1656 => x"30303030",		-- colors: 48, 48, 48, 48
        1657 => x"30303030",		-- colors: 48, 48, 48, 48
        1658 => x"30303032",		-- colors: 48, 48, 48, 50
        1659 => x"30303030",		-- colors: 48, 48, 48, 48
        1660 => x"30303030",		-- colors: 48, 48, 48, 48
        1661 => x"30303030",		-- colors: 48, 48, 48, 48
        1662 => x"30303030",		-- colors: 48, 48, 48, 48

                --  sprite 5
        1663 => x"31313131",		-- colors: 49, 49, 49, 49
        1664 => x"31313030",		-- colors: 49, 49, 48, 48
        1665 => x"30303030",		-- colors: 48, 48, 48, 48
        1666 => x"30303030",		-- colors: 48, 48, 48, 48
        1667 => x"31323131",		-- colors: 49, 50, 49, 49
        1668 => x"31303030",		-- colors: 49, 48, 48, 48
        1669 => x"30303030",		-- colors: 48, 48, 48, 48
        1670 => x"30303030",		-- colors: 48, 48, 48, 48
        1671 => x"32313131",		-- colors: 50, 49, 49, 49
        1672 => x"31303030",		-- colors: 49, 48, 48, 48
        1673 => x"30303030",		-- colors: 48, 48, 48, 48
        1674 => x"30303030",		-- colors: 48, 48, 48, 48
        1675 => x"32313131",		-- colors: 50, 49, 49, 49
        1676 => x"31303030",		-- colors: 49, 48, 48, 48
        1677 => x"30303030",		-- colors: 48, 48, 48, 48
        1678 => x"30303030",		-- colors: 48, 48, 48, 48
        1679 => x"31323131",		-- colors: 49, 50, 49, 49
        1680 => x"32303030",		-- colors: 50, 48, 48, 48
        1681 => x"30303030",		-- colors: 48, 48, 48, 48
        1682 => x"30303030",		-- colors: 48, 48, 48, 48
        1683 => x"32313131",		-- colors: 50, 49, 49, 49
        1684 => x"31323030",		-- colors: 49, 50, 48, 48
        1685 => x"30303030",		-- colors: 48, 48, 48, 48
        1686 => x"30303030",		-- colors: 48, 48, 48, 48
        1687 => x"31313131",		-- colors: 49, 49, 49, 49
        1688 => x"31313230",		-- colors: 49, 49, 50, 48
        1689 => x"30303030",		-- colors: 48, 48, 48, 48
        1690 => x"30303030",		-- colors: 48, 48, 48, 48
        1691 => x"31313131",		-- colors: 49, 49, 49, 49
        1692 => x"31313132",		-- colors: 49, 49, 49, 50
        1693 => x"30303030",		-- colors: 48, 48, 48, 48
        1694 => x"30303030",		-- colors: 48, 48, 48, 48
        1695 => x"31313131",		-- colors: 49, 49, 49, 49
        1696 => x"31313131",		-- colors: 49, 49, 49, 49
        1697 => x"32303030",		-- colors: 50, 48, 48, 48
        1698 => x"30303030",		-- colors: 48, 48, 48, 48
        1699 => x"31313131",		-- colors: 49, 49, 49, 49
        1700 => x"31313131",		-- colors: 49, 49, 49, 49
        1701 => x"32303030",		-- colors: 50, 48, 48, 48
        1702 => x"30303030",		-- colors: 48, 48, 48, 48
        1703 => x"31313131",		-- colors: 49, 49, 49, 49
        1704 => x"31313131",		-- colors: 49, 49, 49, 49
        1705 => x"32303030",		-- colors: 50, 48, 48, 48
        1706 => x"30303030",		-- colors: 48, 48, 48, 48
        1707 => x"31313131",		-- colors: 49, 49, 49, 49
        1708 => x"31313131",		-- colors: 49, 49, 49, 49
        1709 => x"30303030",		-- colors: 48, 48, 48, 48
        1710 => x"30303030",		-- colors: 48, 48, 48, 48
        1711 => x"31313131",		-- colors: 49, 49, 49, 49
        1712 => x"31313131",		-- colors: 49, 49, 49, 49
        1713 => x"30303030",		-- colors: 48, 48, 48, 48
        1714 => x"30303030",		-- colors: 48, 48, 48, 48
        1715 => x"31323231",		-- colors: 49, 50, 50, 49
        1716 => x"31313232",		-- colors: 49, 49, 50, 50
        1717 => x"31323030",		-- colors: 49, 50, 48, 48
        1718 => x"30303030",		-- colors: 48, 48, 48, 48
        1719 => x"32313232",		-- colors: 50, 49, 50, 50
        1720 => x"32323132",		-- colors: 50, 50, 49, 50
        1721 => x"32313230",		-- colors: 50, 49, 50, 48
        1722 => x"30303030",		-- colors: 48, 48, 48, 48
        1723 => x"32323232",		-- colors: 50, 50, 50, 50
        1724 => x"32323232",		-- colors: 50, 50, 50, 50
        1725 => x"32323132",		-- colors: 50, 50, 49, 50
        1726 => x"30303030",		-- colors: 48, 48, 48, 48

				--**mario**

                --  sprite 0
        1727 => x"00000000",		-- colors: 52, 52, 52, 52
        1728 => x"00000000",		-- colors: 52, 52, 52, 52
        1729 => x"00000000",		-- colors: 52, 52, 52, 52
        1730 => x"00000000",		-- colors: 52, 52, 52, 52
        1731 => x"00000000",		-- colors: 52, 52, 52, 52
        1732 => x"00003535",		-- colors: 52, 52, 53, 53
        1733 => x"35350000",		-- colors: 53, 53, 52, 52
        1734 => x"00000000",		-- colors: 52, 52, 52, 52
        1735 => x"00000000",		-- colors: 52, 52, 52, 52
        1736 => x"00353535",		-- colors: 52, 53, 53, 53
        1737 => x"35353535",		-- colors: 53, 53, 53, 53
        1738 => x"35000000",		-- colors: 53, 52, 52, 52
        1739 => x"00000000",		-- colors: 52, 52, 52, 52
        1740 => x"00373737",		-- colors: 52, 55, 55, 55
        1741 => x"37363600",		-- colors: 55, 54, 54, 52
        1742 => x"00000000",		-- colors: 52, 52, 52, 52
        1743 => x"00000000",		-- colors: 52, 52, 52, 52
        1744 => x"37363637",		-- colors: 55, 54, 54, 55
        1745 => x"36363736",		-- colors: 54, 54, 55, 54
        1746 => x"36360000",		-- colors: 54, 54, 52, 52
        1747 => x"00000000",		-- colors: 52, 52, 52, 52
        1748 => x"37363637",		-- colors: 55, 54, 54, 55
        1749 => x"37363637",		-- colors: 55, 54, 54, 55
        1750 => x"36363600",		-- colors: 54, 54, 54, 52
        1751 => x"00000037",		-- colors: 52, 52, 52, 55
        1752 => x"37373636",		-- colors: 55, 55, 54, 54
        1753 => x"36363737",		-- colors: 54, 54, 55, 55
        1754 => x"37370000",		-- colors: 55, 55, 52, 52
        1755 => x"00000000",		-- colors: 52, 52, 52, 52
        1756 => x"00003636",		-- colors: 52, 52, 54, 54
        1757 => x"36363636",		-- colors: 54, 54, 54, 54
        1758 => x"36000000",		-- colors: 54, 52, 52, 52
        1759 => x"00000000",		-- colors: 52, 52, 52, 52
        1760 => x"37373737",		-- colors: 55, 55, 55, 55
        1761 => x"37350036",		-- colors: 55, 53, 52, 54
        1762 => x"00000000",		-- colors: 52, 52, 52, 52
        1763 => x"00000036",		-- colors: 52, 52, 52, 54
        1764 => x"37373737",		-- colors: 55, 55, 55, 55
        1765 => x"37373636",		-- colors: 55, 55, 54, 54
        1766 => x"36000000",		-- colors: 54, 52, 52, 52
        1767 => x"00003636",		-- colors: 52, 52, 54, 54
        1768 => x"35353737",		-- colors: 53, 53, 55, 55
        1769 => x"37373636",		-- colors: 55, 55, 54, 54
        1770 => x"00000000",		-- colors: 52, 52, 52, 52
        1771 => x"37373535",		-- colors: 55, 55, 53, 53
        1772 => x"35353535",		-- colors: 53, 53, 53, 53
        1773 => x"35353535",		-- colors: 53, 53, 53, 53
        1774 => x"00000000",		-- colors: 52, 52, 52, 52
        1775 => x"37373535",		-- colors: 55, 55, 53, 53
        1776 => x"35353535",		-- colors: 53, 53, 53, 53
        1777 => x"35353535",		-- colors: 53, 53, 53, 53
        1778 => x"00000000",		-- colors: 52, 52, 52, 52
        1779 => x"37373535",		-- colors: 55, 55, 53, 53
        1780 => x"35350000",		-- colors: 53, 53, 52, 52
        1781 => x"35353500",		-- colors: 53, 53, 53, 52
        1782 => x"00000000",		-- colors: 52, 52, 52, 52
        1783 => x"37000000",		-- colors: 55, 52, 52, 52
        1784 => x"00000037",		-- colors: 52, 52, 52, 55
        1785 => x"37370000",		-- colors: 55, 55, 52, 52
        1786 => x"00000000",		-- colors: 52, 52, 52, 52
        1787 => x"00000000",		-- colors: 52, 52, 52, 52
        1788 => x"00000037",		-- colors: 52, 52, 52, 55
        1789 => x"37373700",		-- colors: 55, 55, 55, 52
        1790 => x"00000000",		-- colors: 52, 52, 52, 52

                --  sprite 1
        1791 => x"00000000",		-- colors: 52, 52, 52, 52
        1792 => x"00353535",		-- colors: 52, 53, 53, 53
        1793 => x"35000000",		-- colors: 53, 52, 52, 52
        1794 => x"00000000",		-- colors: 52, 52, 52, 52
        1795 => x"00000000",		-- colors: 52, 52, 52, 52
        1796 => x"35353535",		-- colors: 53, 53, 53, 53
        1797 => x"35353535",		-- colors: 53, 53, 53, 53
        1798 => x"00000000",		-- colors: 52, 52, 52, 52
        1799 => x"00000000",		-- colors: 52, 52, 52, 52
        1800 => x"37373737",		-- colors: 55, 55, 55, 55
        1801 => x"36360000",		-- colors: 54, 54, 52, 52
        1802 => x"00000000",		-- colors: 52, 52, 52, 52
        1803 => x"00000037",		-- colors: 52, 52, 52, 55
        1804 => x"36363736",		-- colors: 54, 54, 55, 54
        1805 => x"36373636",		-- colors: 54, 55, 54, 54
        1806 => x"36000000",		-- colors: 54, 52, 52, 52
        1807 => x"00000037",		-- colors: 52, 52, 52, 55
        1808 => x"36363737",		-- colors: 54, 54, 55, 55
        1809 => x"36363736",		-- colors: 54, 54, 55, 54
        1810 => x"36360000",		-- colors: 54, 54, 52, 52
        1811 => x"00003737",		-- colors: 52, 52, 55, 55
        1812 => x"37363636",		-- colors: 55, 54, 54, 54
        1813 => x"36373737",		-- colors: 54, 55, 55, 55
        1814 => x"37000000",		-- colors: 55, 52, 52, 52
        1815 => x"00000000",		-- colors: 52, 52, 52, 52
        1816 => x"00363636",		-- colors: 52, 54, 54, 54
        1817 => x"36363636",		-- colors: 54, 54, 54, 54
        1818 => x"00000000",		-- colors: 52, 52, 52, 52
        1819 => x"00000000",		-- colors: 52, 52, 52, 52
        1820 => x"37373737",		-- colors: 55, 55, 55, 55
        1821 => x"37370000",		-- colors: 55, 55, 52, 52
        1822 => x"00000000",		-- colors: 52, 52, 52, 52
        1823 => x"00000037",		-- colors: 52, 52, 52, 55
        1824 => x"37373735",		-- colors: 55, 55, 55, 53
        1825 => x"35373700",		-- colors: 53, 55, 55, 52
        1826 => x"00000000",		-- colors: 52, 52, 52, 52
        1827 => x"00000037",		-- colors: 52, 52, 52, 55
        1828 => x"37373535",		-- colors: 55, 55, 53, 53
        1829 => x"36353500",		-- colors: 54, 53, 53, 52
        1830 => x"00000000",		-- colors: 52, 52, 52, 52
        1831 => x"00000037",		-- colors: 52, 52, 52, 55
        1832 => x"37373735",		-- colors: 55, 55, 55, 53
        1833 => x"35353535",		-- colors: 53, 53, 53, 53
        1834 => x"00000000",		-- colors: 52, 52, 52, 52
        1835 => x"00000035",		-- colors: 52, 52, 52, 53
        1836 => x"37363636",		-- colors: 55, 54, 54, 54
        1837 => x"35353535",		-- colors: 53, 53, 53, 53
        1838 => x"00000000",		-- colors: 52, 52, 52, 52
        1839 => x"00000035",		-- colors: 52, 52, 52, 53
        1840 => x"35363635",		-- colors: 53, 54, 54, 53
        1841 => x"35353535",		-- colors: 53, 53, 53, 53
        1842 => x"00000000",		-- colors: 52, 52, 52, 52
        1843 => x"00000035",		-- colors: 52, 52, 52, 53
        1844 => x"35353500",		-- colors: 53, 53, 53, 52
        1845 => x"35353500",		-- colors: 53, 53, 53, 52
        1846 => x"00000000",		-- colors: 52, 52, 52, 52
        1847 => x"00000037",		-- colors: 52, 52, 52, 55
        1848 => x"37370000",		-- colors: 55, 55, 52, 52
        1849 => x"37373700",		-- colors: 55, 55, 55, 52
        1850 => x"00000000",		-- colors: 52, 52, 52, 52
        1851 => x"00000037",		-- colors: 52, 52, 52, 55
        1852 => x"37373700",		-- colors: 55, 55, 55, 52
        1853 => x"37373737",		-- colors: 55, 55, 55, 55
        1854 => x"00000000",		-- colors: 52, 52, 52, 52

                --  sprite 2
        1855 => x"00000000",		-- colors: 52, 52, 52, 52
        1856 => x"00353535",		-- colors: 52, 53, 53, 53
        1857 => x"35000000",		-- colors: 53, 52, 52, 52
        1858 => x"00000000",		-- colors: 52, 52, 52, 52
        1859 => x"00000000",		-- colors: 52, 52, 52, 52
        1860 => x"35353535",		-- colors: 53, 53, 53, 53
        1861 => x"35353535",		-- colors: 53, 53, 53, 53
        1862 => x"00000000",		-- colors: 52, 52, 52, 52
        1863 => x"00000000",		-- colors: 52, 52, 52, 52
        1864 => x"37373737",		-- colors: 55, 55, 55, 55
        1865 => x"36360000",		-- colors: 54, 54, 52, 52
        1866 => x"00000000",		-- colors: 52, 52, 52, 52
        1867 => x"00000037",		-- colors: 52, 52, 52, 55
        1868 => x"36363736",		-- colors: 54, 54, 55, 54
        1869 => x"36373636",		-- colors: 54, 55, 54, 54
        1870 => x"36000000",		-- colors: 54, 52, 52, 52
        1871 => x"00000037",		-- colors: 52, 52, 52, 55
        1872 => x"36363737",		-- colors: 54, 54, 55, 55
        1873 => x"36363736",		-- colors: 54, 54, 55, 54
        1874 => x"36360000",		-- colors: 54, 54, 52, 52
        1875 => x"00003737",		-- colors: 52, 52, 55, 55
        1876 => x"37363636",		-- colors: 55, 54, 54, 54
        1877 => x"36373737",		-- colors: 54, 55, 55, 55
        1878 => x"37000000",		-- colors: 55, 52, 52, 52
        1879 => x"00000000",		-- colors: 52, 52, 52, 52
        1880 => x"00363636",		-- colors: 52, 54, 54, 54
        1881 => x"36363636",		-- colors: 54, 54, 54, 54
        1882 => x"00000000",		-- colors: 52, 52, 52, 52
        1883 => x"00003737",		-- colors: 52, 52, 55, 55
        1884 => x"37373535",		-- colors: 55, 55, 53, 53
        1885 => x"37370000",		-- colors: 55, 55, 52, 52
        1886 => x"00363600",		-- colors: 52, 54, 54, 52
        1887 => x"36363737",		-- colors: 54, 54, 55, 55
        1888 => x"37373535",		-- colors: 55, 55, 53, 53
        1889 => x"35373737",		-- colors: 53, 55, 55, 55
        1890 => x"36363600",		-- colors: 54, 54, 54, 52
        1891 => x"36363600",		-- colors: 54, 54, 54, 52
        1892 => x"37373536",		-- colors: 55, 55, 53, 54
        1893 => x"35353537",		-- colors: 53, 53, 53, 55
        1894 => x"37363600",		-- colors: 55, 54, 54, 52
        1895 => x"36360000",		-- colors: 54, 54, 52, 52
        1896 => x"35353535",		-- colors: 53, 53, 53, 53
        1897 => x"35353500",		-- colors: 53, 53, 53, 52
        1898 => x"00370000",		-- colors: 52, 55, 52, 52
        1899 => x"00000035",		-- colors: 52, 52, 52, 53
        1900 => x"35353535",		-- colors: 53, 53, 53, 53
        1901 => x"35353535",		-- colors: 53, 53, 53, 53
        1902 => x"37370000",		-- colors: 55, 55, 52, 52
        1903 => x"00003535",		-- colors: 52, 52, 53, 53
        1904 => x"35353535",		-- colors: 53, 53, 53, 53
        1905 => x"35353535",		-- colors: 53, 53, 53, 53
        1906 => x"37370000",		-- colors: 55, 55, 52, 52
        1907 => x"00373737",		-- colors: 52, 55, 55, 55
        1908 => x"35350000",		-- colors: 53, 53, 52, 52
        1909 => x"00353535",		-- colors: 52, 53, 53, 53
        1910 => x"37370000",		-- colors: 55, 55, 52, 52
        1911 => x"00373737",		-- colors: 52, 55, 55, 55
        1912 => x"00000000",		-- colors: 52, 52, 52, 52
        1913 => x"00000000",		-- colors: 52, 52, 52, 52
        1914 => x"00000000",		-- colors: 52, 52, 52, 52
        1915 => x"00003737",		-- colors: 52, 52, 55, 55
        1916 => x"37000000",		-- colors: 55, 52, 52, 52
        1917 => x"00000000",		-- colors: 52, 52, 52, 52
        1918 => x"00000000",		-- colors: 52, 52, 52, 52

                --  sprite 3
        1919 => x"00000000",		-- colors: 52, 52, 52, 52
        1920 => x"00000000",		-- colors: 52, 52, 52, 52
        1921 => x"00000000",		-- colors: 52, 52, 52, 52
        1922 => x"00000000",		-- colors: 52, 52, 52, 52
        1923 => x"00000000",		-- colors: 52, 52, 52, 52
        1924 => x"00003535",		-- colors: 52, 52, 53, 53
        1925 => x"35350000",		-- colors: 53, 53, 52, 52
        1926 => x"00000000",		-- colors: 52, 52, 52, 52
        1927 => x"00000000",		-- colors: 52, 52, 52, 52
        1928 => x"00353535",		-- colors: 52, 53, 53, 53
        1929 => x"35353535",		-- colors: 53, 53, 53, 53
        1930 => x"35000000",		-- colors: 53, 52, 52, 52
        1931 => x"00000000",		-- colors: 52, 52, 52, 52
        1932 => x"00373737",		-- colors: 52, 55, 55, 55
        1933 => x"37363600",		-- colors: 55, 54, 54, 52
        1934 => x"00000000",		-- colors: 52, 52, 52, 52
        1935 => x"00000000",		-- colors: 52, 52, 52, 52
        1936 => x"37363637",		-- colors: 55, 54, 54, 55
        1937 => x"36363736",		-- colors: 54, 54, 55, 54
        1938 => x"36360000",		-- colors: 54, 54, 52, 52
        1939 => x"00000000",		-- colors: 52, 52, 52, 52
        1940 => x"37363637",		-- colors: 55, 54, 54, 55
        1941 => x"37363637",		-- colors: 55, 54, 54, 55
        1942 => x"36363600",		-- colors: 54, 54, 54, 52
        1943 => x"00000037",		-- colors: 52, 52, 52, 55
        1944 => x"37373636",		-- colors: 55, 55, 54, 54
        1945 => x"36363737",		-- colors: 54, 54, 55, 55
        1946 => x"37370000",		-- colors: 55, 55, 52, 52
        1947 => x"00363600",		-- colors: 52, 54, 54, 52
        1948 => x"00003636",		-- colors: 52, 52, 54, 54
        1949 => x"36363636",		-- colors: 54, 54, 54, 54
        1950 => x"36003636",		-- colors: 54, 52, 54, 54
        1951 => x"36363637",		-- colors: 54, 54, 54, 55
        1952 => x"37373737",		-- colors: 55, 55, 55, 55
        1953 => x"35373700",		-- colors: 53, 55, 55, 52
        1954 => x"00373636",		-- colors: 52, 55, 54, 54
        1955 => x"00003600",		-- colors: 52, 52, 54, 52
        1956 => x"37373735",		-- colors: 55, 55, 55, 53
        1957 => x"35353737",		-- colors: 53, 53, 55, 55
        1958 => x"37373700",		-- colors: 55, 55, 55, 52
        1959 => x"00000000",		-- colors: 52, 52, 52, 52
        1960 => x"00373735",		-- colors: 52, 55, 55, 53
        1961 => x"36353535",		-- colors: 54, 53, 53, 53
        1962 => x"00000000",		-- colors: 52, 52, 52, 52
        1963 => x"00003737",		-- colors: 52, 52, 55, 55
        1964 => x"00353535",		-- colors: 52, 53, 53, 53
        1965 => x"35353535",		-- colors: 53, 53, 53, 53
        1966 => x"00000037",		-- colors: 52, 52, 52, 55
        1967 => x"00373737",		-- colors: 52, 55, 55, 55
        1968 => x"37353535",		-- colors: 55, 53, 53, 53
        1969 => x"35353535",		-- colors: 53, 53, 53, 53
        1970 => x"35353737",		-- colors: 53, 53, 55, 55
        1971 => x"37370035",		-- colors: 55, 55, 52, 53
        1972 => x"35353535",		-- colors: 53, 53, 53, 53
        1973 => x"35353535",		-- colors: 53, 53, 53, 53
        1974 => x"35353737",		-- colors: 53, 53, 55, 55
        1975 => x"00000000",		-- colors: 52, 52, 52, 52
        1976 => x"35353535",		-- colors: 53, 53, 53, 53
        1977 => x"00000000",		-- colors: 52, 52, 52, 52
        1978 => x"00000000",		-- colors: 52, 52, 52, 52
        1979 => x"00000000",		-- colors: 52, 52, 52, 52
        1980 => x"00353500",		-- colors: 52, 53, 53, 52
        1981 => x"00000000",		-- colors: 52, 52, 52, 52
        1982 => x"00000000",		-- colors: 52, 52, 52, 52

                --  sprite 4
        1983 => x"00000000",		-- colors: 52, 52, 52, 52
        1984 => x"00000035",		-- colors: 52, 52, 52, 53
        1985 => x"35353500",		-- colors: 53, 53, 53, 52
        1986 => x"00000000",		-- colors: 52, 52, 52, 52
        1987 => x"00000000",		-- colors: 52, 52, 52, 52
        1988 => x"35353535",		-- colors: 53, 53, 53, 53
        1989 => x"35353535",		-- colors: 53, 53, 53, 53
        1990 => x"00000000",		-- colors: 52, 52, 52, 52
        1991 => x"00000000",		-- colors: 52, 52, 52, 52
        1992 => x"00003636",		-- colors: 52, 52, 54, 54
        1993 => x"37373737",		-- colors: 55, 55, 55, 55
        1994 => x"00000000",		-- colors: 52, 52, 52, 52
        1995 => x"00000036",		-- colors: 52, 52, 52, 54
        1996 => x"36363736",		-- colors: 54, 54, 55, 54
        1997 => x"36373636",		-- colors: 54, 55, 54, 54
        1998 => x"37000000",		-- colors: 55, 52, 52, 52
        1999 => x"00003636",		-- colors: 52, 52, 54, 54
        2000 => x"36373636",		-- colors: 54, 55, 54, 54
        2001 => x"37373636",		-- colors: 55, 55, 54, 54
        2002 => x"37000000",		-- colors: 55, 52, 52, 52
        2003 => x"00000037",		-- colors: 52, 52, 52, 55
        2004 => x"37373736",		-- colors: 55, 55, 55, 54
        2005 => x"36363637",		-- colors: 54, 54, 54, 55
        2006 => x"37370000",		-- colors: 55, 55, 52, 52
        2007 => x"00000000",		-- colors: 52, 52, 52, 52
        2008 => x"36363636",		-- colors: 54, 54, 54, 54
        2009 => x"36363600",		-- colors: 54, 54, 54, 52
        2010 => x"00000000",		-- colors: 52, 52, 52, 52
        2011 => x"00363600",		-- colors: 52, 54, 54, 52
        2012 => x"00003737",		-- colors: 52, 52, 55, 55
        2013 => x"35353737",		-- colors: 53, 53, 55, 55
        2014 => x"37370000",		-- colors: 55, 55, 52, 52
        2015 => x"00363636",		-- colors: 52, 54, 54, 54
        2016 => x"37373735",		-- colors: 55, 55, 55, 53
        2017 => x"35353737",		-- colors: 53, 53, 55, 55
        2018 => x"37373636",		-- colors: 55, 55, 54, 54
        2019 => x"00363637",		-- colors: 52, 54, 54, 55
        2020 => x"37353535",		-- colors: 55, 53, 53, 53
        2021 => x"36353737",		-- colors: 54, 53, 55, 55
        2022 => x"00363636",		-- colors: 52, 54, 54, 54
        2023 => x"00003700",		-- colors: 52, 52, 55, 52
        2024 => x"00353535",		-- colors: 52, 53, 53, 53
        2025 => x"35353535",		-- colors: 53, 53, 53, 53
        2026 => x"00003636",		-- colors: 52, 52, 54, 54
        2027 => x"00003737",		-- colors: 52, 52, 55, 55
        2028 => x"35353535",		-- colors: 53, 53, 53, 53
        2029 => x"35353535",		-- colors: 53, 53, 53, 53
        2030 => x"35000000",		-- colors: 53, 52, 52, 52
        2031 => x"00003737",		-- colors: 52, 52, 55, 55
        2032 => x"35353535",		-- colors: 53, 53, 53, 53
        2033 => x"35353535",		-- colors: 53, 53, 53, 53
        2034 => x"35350000",		-- colors: 53, 53, 52, 52
        2035 => x"00003737",		-- colors: 52, 52, 55, 55
        2036 => x"35353500",		-- colors: 53, 53, 53, 52
        2037 => x"00003535",		-- colors: 52, 52, 53, 53
        2038 => x"37373700",		-- colors: 55, 55, 55, 52
        2039 => x"00000000",		-- colors: 52, 52, 52, 52
        2040 => x"00000000",		-- colors: 52, 52, 52, 52
        2041 => x"00000000",		-- colors: 52, 52, 52, 52
        2042 => x"37373700",		-- colors: 55, 55, 55, 52
        2043 => x"00000000",		-- colors: 52, 52, 52, 52
        2044 => x"00000000",		-- colors: 52, 52, 52, 52
        2045 => x"00000037",		-- colors: 52, 52, 52, 55
        2046 => x"37370000",		-- colors: 55, 55, 52, 52

                --  sprite 5
        2047 => x"00000000",		-- colors: 52, 52, 52, 52
        2048 => x"00000035",		-- colors: 52, 52, 52, 53
        2049 => x"35353500",		-- colors: 53, 53, 53, 52
        2050 => x"00000000",		-- colors: 52, 52, 52, 52
        2051 => x"00000000",		-- colors: 52, 52, 52, 52
        2052 => x"35353535",		-- colors: 53, 53, 53, 53
        2053 => x"35353535",		-- colors: 53, 53, 53, 53
        2054 => x"00000000",		-- colors: 52, 52, 52, 52
        2055 => x"00000000",		-- colors: 52, 52, 52, 52
        2056 => x"00003636",		-- colors: 52, 52, 54, 54
        2057 => x"37373737",		-- colors: 55, 55, 55, 55
        2058 => x"00000000",		-- colors: 52, 52, 52, 52
        2059 => x"00000036",		-- colors: 52, 52, 52, 54
        2060 => x"36363736",		-- colors: 54, 54, 55, 54
        2061 => x"36373636",		-- colors: 54, 55, 54, 54
        2062 => x"37000000",		-- colors: 55, 52, 52, 52
        2063 => x"00003636",		-- colors: 52, 52, 54, 54
        2064 => x"36373636",		-- colors: 54, 55, 54, 54
        2065 => x"37373636",		-- colors: 55, 55, 54, 54
        2066 => x"37000000",		-- colors: 55, 52, 52, 52
        2067 => x"00000037",		-- colors: 52, 52, 52, 55
        2068 => x"37373736",		-- colors: 55, 55, 55, 54
        2069 => x"36363637",		-- colors: 54, 54, 54, 55
        2070 => x"37370000",		-- colors: 55, 55, 52, 52
        2071 => x"00000000",		-- colors: 52, 52, 52, 52
        2072 => x"36363636",		-- colors: 54, 54, 54, 54
        2073 => x"36363600",		-- colors: 54, 54, 54, 52
        2074 => x"00000000",		-- colors: 52, 52, 52, 52
        2075 => x"00000000",		-- colors: 52, 52, 52, 52
        2076 => x"00003737",		-- colors: 52, 52, 55, 55
        2077 => x"37373737",		-- colors: 55, 55, 55, 55
        2078 => x"00000000",		-- colors: 52, 52, 52, 52
        2079 => x"00000000",		-- colors: 52, 52, 52, 52
        2080 => x"00373735",		-- colors: 52, 55, 55, 53
        2081 => x"35373737",		-- colors: 53, 55, 55, 55
        2082 => x"37000000",		-- colors: 55, 52, 52, 52
        2083 => x"00000000",		-- colors: 52, 52, 52, 52
        2084 => x"00353536",		-- colors: 52, 53, 53, 54
        2085 => x"35353737",		-- colors: 53, 53, 55, 55
        2086 => x"37000000",		-- colors: 55, 52, 52, 52
        2087 => x"00000000",		-- colors: 52, 52, 52, 52
        2088 => x"35353535",		-- colors: 53, 53, 53, 53
        2089 => x"35373737",		-- colors: 53, 55, 55, 55
        2090 => x"37000000",		-- colors: 55, 52, 52, 52
        2091 => x"00000000",		-- colors: 52, 52, 52, 52
        2092 => x"35353535",		-- colors: 53, 53, 53, 53
        2093 => x"36363637",		-- colors: 54, 54, 54, 55
        2094 => x"35000000",		-- colors: 53, 52, 52, 52
        2095 => x"00000000",		-- colors: 52, 52, 52, 52
        2096 => x"35353535",		-- colors: 53, 53, 53, 53
        2097 => x"35363635",		-- colors: 53, 54, 54, 53
        2098 => x"35000000",		-- colors: 53, 52, 52, 52
        2099 => x"00000000",		-- colors: 52, 52, 52, 52
        2100 => x"00353535",		-- colors: 52, 53, 53, 53
        2101 => x"00353535",		-- colors: 52, 53, 53, 53
        2102 => x"35000000",		-- colors: 53, 52, 52, 52
        2103 => x"00000000",		-- colors: 52, 52, 52, 52
        2104 => x"00373737",		-- colors: 52, 55, 55, 55
        2105 => x"00003737",		-- colors: 52, 52, 55, 55
        2106 => x"37000000",		-- colors: 55, 52, 52, 52
        2107 => x"00000000",		-- colors: 52, 52, 52, 52
        2108 => x"37373737",		-- colors: 55, 55, 55, 55
        2109 => x"00373737",		-- colors: 52, 55, 55, 55
        2110 => x"37000000",		-- colors: 55, 52, 52, 52

                --  sprite 6
        2111 => x"00000000",		-- colors: 52, 52, 52, 52
        2112 => x"00000000",		-- colors: 52, 52, 52, 52
        2113 => x"00000000",		-- colors: 52, 52, 52, 52
        2114 => x"00000000",		-- colors: 52, 52, 52, 52
        2115 => x"00000000",		-- colors: 52, 52, 52, 52
        2116 => x"00003535",		-- colors: 52, 52, 53, 53
        2117 => x"35350000",		-- colors: 53, 53, 52, 52
        2118 => x"00000000",		-- colors: 52, 52, 52, 52
        2119 => x"00000035",		-- colors: 52, 52, 52, 53
        2120 => x"35353535",		-- colors: 53, 53, 53, 53
        2121 => x"35353500",		-- colors: 53, 53, 53, 52
        2122 => x"00000000",		-- colors: 52, 52, 52, 52
        2123 => x"00000000",		-- colors: 52, 52, 52, 52
        2124 => x"00363637",		-- colors: 52, 54, 54, 55
        2125 => x"37373700",		-- colors: 55, 55, 55, 52
        2126 => x"00000000",		-- colors: 52, 52, 52, 52
        2127 => x"00003636",		-- colors: 52, 52, 54, 54
        2128 => x"36373636",		-- colors: 54, 55, 54, 54
        2129 => x"37363637",		-- colors: 55, 54, 54, 55
        2130 => x"00000000",		-- colors: 52, 52, 52, 52
        2131 => x"00363636",		-- colors: 52, 54, 54, 54
        2132 => x"37363637",		-- colors: 55, 54, 54, 55
        2133 => x"37363637",		-- colors: 55, 54, 54, 55
        2134 => x"00000000",		-- colors: 52, 52, 52, 52
        2135 => x"00003737",		-- colors: 52, 52, 55, 55
        2136 => x"37373636",		-- colors: 55, 55, 54, 54
        2137 => x"36363737",		-- colors: 54, 54, 55, 55
        2138 => x"37000000",		-- colors: 55, 52, 52, 52
        2139 => x"00000036",		-- colors: 52, 52, 52, 54
        2140 => x"36363636",		-- colors: 54, 54, 54, 54
        2141 => x"36360000",		-- colors: 54, 54, 52, 52
        2142 => x"00000000",		-- colors: 52, 52, 52, 52
        2143 => x"00000000",		-- colors: 52, 52, 52, 52
        2144 => x"36003537",		-- colors: 54, 52, 53, 55
        2145 => x"37373737",		-- colors: 55, 55, 55, 55
        2146 => x"00000000",		-- colors: 52, 52, 52, 52
        2147 => x"00000036",		-- colors: 52, 52, 52, 54
        2148 => x"36363737",		-- colors: 54, 54, 55, 55
        2149 => x"37373737",		-- colors: 55, 55, 55, 55
        2150 => x"36000000",		-- colors: 54, 52, 52, 52
        2151 => x"00000000",		-- colors: 52, 52, 52, 52
        2152 => x"36363737",		-- colors: 54, 54, 55, 55
        2153 => x"37373535",		-- colors: 55, 55, 53, 53
        2154 => x"36360000",		-- colors: 54, 54, 52, 52
        2155 => x"00000000",		-- colors: 52, 52, 52, 52
        2156 => x"35353535",		-- colors: 53, 53, 53, 53
        2157 => x"35353535",		-- colors: 53, 53, 53, 53
        2158 => x"35353737",		-- colors: 53, 53, 55, 55
        2159 => x"00000000",		-- colors: 52, 52, 52, 52
        2160 => x"35353535",		-- colors: 53, 53, 53, 53
        2161 => x"35353535",		-- colors: 53, 53, 53, 53
        2162 => x"35353737",		-- colors: 53, 53, 55, 55
        2163 => x"00000000",		-- colors: 52, 52, 52, 52
        2164 => x"00353535",		-- colors: 52, 53, 53, 53
        2165 => x"00003535",		-- colors: 52, 52, 53, 53
        2166 => x"35353737",		-- colors: 53, 53, 55, 55
        2167 => x"00000000",		-- colors: 52, 52, 52, 52
        2168 => x"00003737",		-- colors: 52, 52, 55, 55
        2169 => x"37000000",		-- colors: 55, 52, 52, 52
        2170 => x"00000037",		-- colors: 52, 52, 52, 55
        2171 => x"00000000",		-- colors: 52, 52, 52, 52
        2172 => x"00373737",		-- colors: 52, 55, 55, 55
        2173 => x"37000000",		-- colors: 55, 52, 52, 52
        2174 => x"00000000",		-- colors: 52, 52, 52, 52

                --  sprite 7
        2175 => x"00000000",		-- colors: 52, 52, 52, 52
        2176 => x"00000000",		-- colors: 52, 52, 52, 52
        2177 => x"00000000",		-- colors: 52, 52, 52, 52
        2178 => x"00000000",		-- colors: 52, 52, 52, 52
        2179 => x"00000000",		-- colors: 52, 52, 52, 52
        2180 => x"00003535",		-- colors: 52, 52, 53, 53
        2181 => x"35350000",		-- colors: 53, 53, 52, 52
        2182 => x"00000000",		-- colors: 52, 52, 52, 52
        2183 => x"00000035",		-- colors: 52, 52, 52, 53
        2184 => x"35353535",		-- colors: 53, 53, 53, 53
        2185 => x"35353500",		-- colors: 53, 53, 53, 52
        2186 => x"00000000",		-- colors: 52, 52, 52, 52
        2187 => x"00000000",		-- colors: 52, 52, 52, 52
        2188 => x"00363637",		-- colors: 52, 54, 54, 55
        2189 => x"37373700",		-- colors: 55, 55, 55, 52
        2190 => x"00000000",		-- colors: 52, 52, 52, 52
        2191 => x"00003636",		-- colors: 52, 52, 54, 54
        2192 => x"36373636",		-- colors: 54, 55, 54, 54
        2193 => x"37363637",		-- colors: 55, 54, 54, 55
        2194 => x"00000000",		-- colors: 52, 52, 52, 52
        2195 => x"00363636",		-- colors: 52, 54, 54, 54
        2196 => x"37363637",		-- colors: 55, 54, 54, 55
        2197 => x"37363637",		-- colors: 55, 54, 54, 55
        2198 => x"00000000",		-- colors: 52, 52, 52, 52
        2199 => x"00003737",		-- colors: 52, 52, 55, 55
        2200 => x"37373636",		-- colors: 55, 55, 54, 54
        2201 => x"36363737",		-- colors: 54, 54, 55, 55
        2202 => x"37000000",		-- colors: 55, 52, 52, 52
        2203 => x"36360036",		-- colors: 54, 54, 52, 54
        2204 => x"36363636",		-- colors: 54, 54, 54, 54
        2205 => x"36360000",		-- colors: 54, 54, 52, 52
        2206 => x"00363600",		-- colors: 52, 54, 54, 52
        2207 => x"36363700",		-- colors: 54, 54, 55, 52
        2208 => x"00373735",		-- colors: 52, 55, 55, 53
        2209 => x"37373737",		-- colors: 55, 55, 55, 55
        2210 => x"37363636",		-- colors: 55, 54, 54, 54
        2211 => x"00373737",		-- colors: 52, 55, 55, 55
        2212 => x"37373535",		-- colors: 55, 55, 53, 53
        2213 => x"35373737",		-- colors: 53, 55, 55, 55
        2214 => x"00360000",		-- colors: 52, 54, 52, 52
        2215 => x"00000000",		-- colors: 52, 52, 52, 52
        2216 => x"35353536",		-- colors: 53, 53, 53, 54
        2217 => x"35373700",		-- colors: 53, 55, 55, 52
        2218 => x"00000000",		-- colors: 52, 52, 52, 52
        2219 => x"37000000",		-- colors: 55, 52, 52, 52
        2220 => x"35353535",		-- colors: 53, 53, 53, 53
        2221 => x"35353500",		-- colors: 53, 53, 53, 52
        2222 => x"37370000",		-- colors: 55, 55, 52, 52
        2223 => x"37373535",		-- colors: 55, 55, 53, 53
        2224 => x"35353535",		-- colors: 53, 53, 53, 53
        2225 => x"35353537",		-- colors: 53, 53, 53, 55
        2226 => x"37373700",		-- colors: 55, 55, 55, 52
        2227 => x"37373535",		-- colors: 55, 55, 53, 53
        2228 => x"35353535",		-- colors: 53, 53, 53, 53
        2229 => x"35353535",		-- colors: 53, 53, 53, 53
        2230 => x"35003737",		-- colors: 53, 52, 55, 55
        2231 => x"00000000",		-- colors: 52, 52, 52, 52
        2232 => x"00000000",		-- colors: 52, 52, 52, 52
        2233 => x"35353535",		-- colors: 53, 53, 53, 53
        2234 => x"00000000",		-- colors: 52, 52, 52, 52
        2235 => x"00000000",		-- colors: 52, 52, 52, 52
        2236 => x"00000000",		-- colors: 52, 52, 52, 52
        2237 => x"00353500",		-- colors: 52, 53, 53, 52
        2238 => x"00000000",		-- colors: 52, 52, 52, 52

                --  sprite 8
        2239 => x"00000000",		-- colors: 52, 52, 52, 52
        2240 => x"00000000",		-- colors: 52, 52, 52, 52
        2241 => x"00000000",		-- colors: 52, 52, 52, 52
        2242 => x"00000000",		-- colors: 52, 52, 52, 52
        2243 => x"00000000",		-- colors: 52, 52, 52, 52
        2244 => x"36363636",		-- colors: 54, 54, 54, 54
        2245 => x"36373700",		-- colors: 54, 55, 55, 52
        2246 => x"00000000",		-- colors: 52, 52, 52, 52
        2247 => x"00003637",		-- colors: 52, 52, 54, 55
        2248 => x"35373737",		-- colors: 53, 55, 55, 55
        2249 => x"37353737",		-- colors: 55, 53, 55, 55
        2250 => x"00000000",		-- colors: 52, 52, 52, 52
        2251 => x"00363735",		-- colors: 52, 54, 55, 53
        2252 => x"35353737",		-- colors: 53, 53, 55, 55
        2253 => x"35353737",		-- colors: 53, 53, 55, 55
        2254 => x"37360000",		-- colors: 55, 54, 52, 52
        2255 => x"00003535",		-- colors: 52, 52, 53, 53
        2256 => x"35353535",		-- colors: 53, 53, 53, 53
        2257 => x"35353535",		-- colors: 53, 53, 53, 53
        2258 => x"37363600",		-- colors: 55, 54, 54, 52
        2259 => x"00353535",		-- colors: 52, 53, 53, 53
        2260 => x"35353535",		-- colors: 53, 53, 53, 53
        2261 => x"35353535",		-- colors: 53, 53, 53, 53
        2262 => x"35363600",		-- colors: 53, 54, 54, 52
        2263 => x"00353535",		-- colors: 52, 53, 53, 53
        2264 => x"35353535",		-- colors: 53, 53, 53, 53
        2265 => x"35353535",		-- colors: 53, 53, 53, 53
        2266 => x"35350000",		-- colors: 53, 53, 52, 52
        2267 => x"00353535",		-- colors: 52, 53, 53, 53
        2268 => x"35353535",		-- colors: 53, 53, 53, 53
        2269 => x"35353535",		-- colors: 53, 53, 53, 53
        2270 => x"35350000",		-- colors: 53, 53, 52, 52
        2271 => x"00353535",		-- colors: 52, 53, 53, 53
        2272 => x"35353535",		-- colors: 53, 53, 53, 53
        2273 => x"35353535",		-- colors: 53, 53, 53, 53
        2274 => x"35000000",		-- colors: 53, 52, 52, 52
        2275 => x"00003535",		-- colors: 52, 52, 53, 53
        2276 => x"35353500",		-- colors: 53, 53, 53, 52
        2277 => x"35353535",		-- colors: 53, 53, 53, 53
        2278 => x"00000000",		-- colors: 52, 52, 52, 52
        2279 => x"00000035",		-- colors: 52, 52, 52, 53
        2280 => x"35353535",		-- colors: 53, 53, 53, 53
        2281 => x"37373737",		-- colors: 55, 55, 55, 55
        2282 => x"00000000",		-- colors: 52, 52, 52, 52
        2283 => x"00000035",		-- colors: 52, 52, 52, 53
        2284 => x"35353535",		-- colors: 53, 53, 53, 53
        2285 => x"37373700",		-- colors: 55, 55, 55, 52
        2286 => x"00000000",		-- colors: 52, 52, 52, 52
        2287 => x"00000000",		-- colors: 52, 52, 52, 52
        2288 => x"35373737",		-- colors: 53, 55, 55, 55
        2289 => x"35000000",		-- colors: 53, 52, 52, 52
        2290 => x"00000000",		-- colors: 52, 52, 52, 52
        2291 => x"00000000",		-- colors: 52, 52, 52, 52
        2292 => x"37373737",		-- colors: 55, 55, 55, 55
        2293 => x"37000000",		-- colors: 55, 52, 52, 52
        2294 => x"00000000",		-- colors: 52, 52, 52, 52
        2295 => x"00000000",		-- colors: 52, 52, 52, 52
        2296 => x"37373737",		-- colors: 55, 55, 55, 55
        2297 => x"37370000",		-- colors: 55, 55, 52, 52
        2298 => x"00000000",		-- colors: 52, 52, 52, 52
        2299 => x"00000000",		-- colors: 52, 52, 52, 52
        2300 => x"00373737",		-- colors: 52, 55, 55, 55
        2301 => x"37370000",		-- colors: 55, 55, 52, 52
        2302 => x"00000000",		-- colors: 52, 52, 52, 52

                --  sprite 9
        2303 => x"00000000",		-- colors: 52, 52, 52, 52
        2304 => x"00000000",		-- colors: 52, 52, 52, 52
        2305 => x"00000000",		-- colors: 52, 52, 52, 52
        2306 => x"00000000",		-- colors: 52, 52, 52, 52
        2307 => x"00000000",		-- colors: 52, 52, 52, 52
        2308 => x"00353535",		-- colors: 52, 53, 53, 53
        2309 => x"35353500",		-- colors: 53, 53, 53, 52
        2310 => x"00000000",		-- colors: 52, 52, 52, 52
        2311 => x"00000000",		-- colors: 52, 52, 52, 52
        2312 => x"00373535",		-- colors: 52, 55, 53, 53
        2313 => x"35353700",		-- colors: 53, 53, 55, 52
        2314 => x"00000000",		-- colors: 52, 52, 52, 52
        2315 => x"00000000",		-- colors: 52, 52, 52, 52
        2316 => x"37373737",		-- colors: 55, 55, 55, 55
        2317 => x"37373737",		-- colors: 55, 55, 55, 55
        2318 => x"00000000",		-- colors: 52, 52, 52, 52
        2319 => x"00000000",		-- colors: 52, 52, 52, 52
        2320 => x"37373737",		-- colors: 55, 55, 55, 55
        2321 => x"37373737",		-- colors: 55, 55, 55, 55
        2322 => x"00000000",		-- colors: 52, 52, 52, 52
        2323 => x"00000000",		-- colors: 52, 52, 52, 52
        2324 => x"00363636",		-- colors: 52, 54, 54, 54
        2325 => x"36363600",		-- colors: 54, 54, 54, 52
        2326 => x"00000000",		-- colors: 52, 52, 52, 52
        2327 => x"00000037",		-- colors: 52, 52, 52, 55
        2328 => x"37353737",		-- colors: 55, 53, 55, 55
        2329 => x"37373537",		-- colors: 55, 55, 53, 55
        2330 => x"37000000",		-- colors: 55, 52, 52, 52
        2331 => x"00003737",		-- colors: 52, 52, 55, 55
        2332 => x"37353737",		-- colors: 55, 53, 55, 55
        2333 => x"37373537",		-- colors: 55, 55, 53, 55
        2334 => x"37370000",		-- colors: 55, 55, 52, 52
        2335 => x"00373737",		-- colors: 52, 55, 55, 55
        2336 => x"35353737",		-- colors: 53, 53, 55, 55
        2337 => x"37373535",		-- colors: 55, 55, 53, 53
        2338 => x"37373700",		-- colors: 55, 55, 55, 52
        2339 => x"36373735",		-- colors: 54, 55, 55, 53
        2340 => x"35353537",		-- colors: 53, 53, 53, 55
        2341 => x"37353535",		-- colors: 55, 53, 53, 53
        2342 => x"35373736",		-- colors: 53, 55, 55, 54
        2343 => x"36363635",		-- colors: 54, 54, 54, 53
        2344 => x"35353535",		-- colors: 53, 53, 53, 53
        2345 => x"35353535",		-- colors: 53, 53, 53, 53
        2346 => x"35363636",		-- colors: 53, 54, 54, 54
        2347 => x"00000035",		-- colors: 52, 52, 52, 53
        2348 => x"35353535",		-- colors: 53, 53, 53, 53
        2349 => x"35353535",		-- colors: 53, 53, 53, 53
        2350 => x"35000000",		-- colors: 53, 52, 52, 52
        2351 => x"00000035",		-- colors: 52, 52, 52, 53
        2352 => x"35353535",		-- colors: 53, 53, 53, 53
        2353 => x"35353535",		-- colors: 53, 53, 53, 53
        2354 => x"35000000",		-- colors: 53, 52, 52, 52
        2355 => x"00000035",		-- colors: 52, 52, 52, 53
        2356 => x"35353500",		-- colors: 53, 53, 53, 52
        2357 => x"00353535",		-- colors: 52, 53, 53, 53
        2358 => x"35000000",		-- colors: 53, 52, 52, 52
        2359 => x"00000000",		-- colors: 52, 52, 52, 52
        2360 => x"35353535",		-- colors: 53, 53, 53, 53
        2361 => x"35353535",		-- colors: 53, 53, 53, 53
        2362 => x"00000000",		-- colors: 52, 52, 52, 52
        2363 => x"00000037",		-- colors: 52, 52, 52, 55
        2364 => x"37373737",		-- colors: 55, 55, 55, 55
        2365 => x"37373737",		-- colors: 55, 55, 55, 55
        2366 => x"37000000",		-- colors: 55, 52, 52, 52


--**princeza**

--  sprite 0
        2367 => x"38383838",		-- colors: 56, 56, 56, 56
        2368 => x"38383939",		-- colors: 56, 56, 57, 57
        2369 => x"39393939",		-- colors: 57, 57, 57, 57
        2370 => x"38383838",		-- colors: 56, 56, 56, 56
        2371 => x"38383838",		-- colors: 56, 56, 56, 56
        2372 => x"38393939",		-- colors: 56, 57, 57, 57
        2373 => x"39393939",		-- colors: 57, 57, 57, 57
        2374 => x"39383838",		-- colors: 57, 56, 56, 56
        2375 => x"39383839",		-- colors: 57, 56, 56, 57
        2376 => x"38393A39",		-- colors: 56, 57, 58, 57
        2377 => x"3A3A3A3A",		-- colors: 58, 58, 58, 58
        2378 => x"38383838",		-- colors: 56, 56, 56, 56
        2379 => x"38393939",		-- colors: 56, 57, 57, 57
        2380 => x"3939393A",		-- colors: 57, 57, 57, 58
        2381 => x"3A3A393A",		-- colors: 58, 58, 57, 58
        2382 => x"3A383838",		-- colors: 58, 56, 56, 56
        2383 => x"38383839",		-- colors: 56, 56, 56, 57
        2384 => x"39393A3A",		-- colors: 57, 57, 58, 58
        2385 => x"3A3A3A3A",		-- colors: 58, 58, 58, 58
        2386 => x"38383838",		-- colors: 56, 56, 56, 56
        2387 => x"38383939",		-- colors: 56, 56, 57, 57
        2388 => x"3938393A",		-- colors: 57, 56, 57, 58
        2389 => x"3A3A3A38",		-- colors: 58, 58, 58, 56
        2390 => x"38383838",		-- colors: 56, 56, 56, 56
        2391 => x"38383838",		-- colors: 56, 56, 56, 56
        2392 => x"38383B3A",		-- colors: 56, 56, 59, 58
        2393 => x"3A383838",		-- colors: 58, 56, 56, 56
        2394 => x"38383838",		-- colors: 56, 56, 56, 56
        2395 => x"38383838",		-- colors: 56, 56, 56, 56
        2396 => x"383B3B3B",		-- colors: 56, 59, 59, 59
        2397 => x"3B383838",		-- colors: 59, 56, 56, 56
        2398 => x"38383838",		-- colors: 56, 56, 56, 56
        2399 => x"38383838",		-- colors: 56, 56, 56, 56
        2400 => x"383B3A3B",		-- colors: 56, 59, 58, 59
        2401 => x"3B3A3838",		-- colors: 59, 58, 56, 56
        2402 => x"38383838",		-- colors: 56, 56, 56, 56
        2403 => x"38383838",		-- colors: 56, 56, 56, 56
        2404 => x"3B3B3B3B",		-- colors: 59, 59, 59, 59
        2405 => x"3B3B3B38",		-- colors: 59, 59, 59, 56
        2406 => x"38383838",		-- colors: 56, 56, 56, 56
        2407 => x"38383838",		-- colors: 56, 56, 56, 56
        2408 => x"3B3B3A3B",		-- colors: 59, 59, 58, 59
        2409 => x"3B3B3B38",		-- colors: 59, 59, 59, 56
        2410 => x"38383838",		-- colors: 56, 56, 56, 56
        2411 => x"3838383B",		-- colors: 56, 56, 56, 59
        2412 => x"3B3A3A3A",		-- colors: 59, 58, 58, 58
        2413 => x"3B3A3A3B",		-- colors: 59, 58, 58, 59
        2414 => x"38383838",		-- colors: 56, 56, 56, 56
        2415 => x"38383B3B",		-- colors: 56, 56, 59, 59
        2416 => x"3B3A3A3B",		-- colors: 59, 58, 58, 59
        2417 => x"3B3B3B3B",		-- colors: 59, 59, 59, 59
        2418 => x"3A383838",		-- colors: 58, 56, 56, 56
        2419 => x"38383A3A",		-- colors: 56, 56, 58, 58
        2420 => x"3B3B3B3B",		-- colors: 59, 59, 59, 59
        2421 => x"3B3A3A3A",		-- colors: 59, 58, 58, 58
        2422 => x"38383838",		-- colors: 56, 56, 56, 56
        2423 => x"38383838",		-- colors: 56, 56, 56, 56
        2424 => x"39393838",		-- colors: 57, 57, 56, 56
        2425 => x"38393938",		-- colors: 56, 57, 57, 56
        2426 => x"38383838",		-- colors: 56, 56, 56, 56
        2427 => x"38383838",		-- colors: 56, 56, 56, 56
        2428 => x"39393938",		-- colors: 57, 57, 57, 56
        2429 => x"38393939",		-- colors: 56, 57, 57, 57
        2430 => x"38383838",		-- colors: 56, 56, 56, 56

                --  sprite 1
        2431 => x"38383838",		-- colors: 56, 56, 56, 56
        2432 => x"38383939",		-- colors: 56, 56, 57, 57
        2433 => x"39393939",		-- colors: 57, 57, 57, 57
        2434 => x"38383838",		-- colors: 56, 56, 56, 56
        2435 => x"38383838",		-- colors: 56, 56, 56, 56
        2436 => x"38393939",		-- colors: 56, 57, 57, 57
        2437 => x"39393939",		-- colors: 57, 57, 57, 57
        2438 => x"39383838",		-- colors: 57, 56, 56, 56
        2439 => x"38383839",		-- colors: 56, 56, 56, 57
        2440 => x"38393A39",		-- colors: 56, 57, 58, 57
        2441 => x"3A3A3A3A",		-- colors: 58, 58, 58, 58
        2442 => x"38383838",		-- colors: 56, 56, 56, 56
        2443 => x"38393939",		-- colors: 56, 57, 57, 57
        2444 => x"3939393A",		-- colors: 57, 57, 57, 58
        2445 => x"3A3A393A",		-- colors: 58, 58, 57, 58
        2446 => x"3A383838",		-- colors: 58, 56, 56, 56
        2447 => x"38383839",		-- colors: 56, 56, 56, 57
        2448 => x"39393A3A",		-- colors: 57, 57, 58, 58
        2449 => x"3A3A3A3A",		-- colors: 58, 58, 58, 58
        2450 => x"38383838",		-- colors: 56, 56, 56, 56
        2451 => x"38393939",		-- colors: 56, 57, 57, 57
        2452 => x"3838393A",		-- colors: 56, 56, 57, 58
        2453 => x"3A3A3A38",		-- colors: 58, 58, 58, 56
        2454 => x"38383838",		-- colors: 56, 56, 56, 56
        2455 => x"38383838",		-- colors: 56, 56, 56, 56
        2456 => x"383B3B3A",		-- colors: 56, 59, 59, 58
        2457 => x"3A383838",		-- colors: 58, 56, 56, 56
        2458 => x"38383838",		-- colors: 56, 56, 56, 56
        2459 => x"3838383B",		-- colors: 56, 56, 56, 59
        2460 => x"3B3B3B3B",		-- colors: 59, 59, 59, 59
        2461 => x"3B3B3838",		-- colors: 59, 59, 56, 56
        2462 => x"3A3A3838",		-- colors: 58, 58, 56, 56
        2463 => x"3A3A3A3B",		-- colors: 58, 58, 58, 59
        2464 => x"3B3B3B3B",		-- colors: 59, 59, 59, 59
        2465 => x"3B3B3B3B",		-- colors: 59, 59, 59, 59
        2466 => x"3A3A3838",		-- colors: 58, 58, 56, 56
        2467 => x"383A3A38",		-- colors: 56, 58, 58, 56
        2468 => x"383B3B3B",		-- colors: 56, 59, 59, 59
        2469 => x"3B3B3B3B",		-- colors: 59, 59, 59, 59
        2470 => x"38383838",		-- colors: 56, 56, 56, 56
        2471 => x"38383838",		-- colors: 56, 56, 56, 56
        2472 => x"3B3B3A3A",		-- colors: 59, 59, 58, 58
        2473 => x"3B3B3B3A",		-- colors: 59, 59, 59, 58
        2474 => x"38393938",		-- colors: 56, 57, 57, 56
        2475 => x"3838383A",		-- colors: 56, 56, 56, 58
        2476 => x"3A3B3B3B",		-- colors: 58, 59, 59, 59
        2477 => x"3B3B3B3B",		-- colors: 59, 59, 59, 59
        2478 => x"39393938",		-- colors: 57, 57, 57, 56
        2479 => x"38383B3B",		-- colors: 56, 56, 59, 59
        2480 => x"3B3B3B3A",		-- colors: 59, 59, 59, 58
        2481 => x"3A3A3A3A",		-- colors: 58, 58, 58, 58
        2482 => x"39393838",		-- colors: 57, 57, 56, 56
        2483 => x"38383A3A",		-- colors: 56, 56, 58, 58
        2484 => x"3A3A3A38",		-- colors: 58, 58, 58, 56
        2485 => x"38383838",		-- colors: 56, 56, 56, 56
        2486 => x"38383838",		-- colors: 56, 56, 56, 56
        2487 => x"38383939",		-- colors: 56, 56, 57, 57
        2488 => x"38383838",		-- colors: 56, 56, 56, 56
        2489 => x"38383838",		-- colors: 56, 56, 56, 56
        2490 => x"38383838",		-- colors: 56, 56, 56, 56
        2491 => x"38383939",		-- colors: 56, 56, 57, 57
        2492 => x"39383838",		-- colors: 57, 56, 56, 56
        2493 => x"38383838",		-- colors: 56, 56, 56, 56
        2494 => x"38383838",		-- colors: 56, 56, 56, 56

                --  sprite 2
        2495 => x"38383838",		-- colors: 56, 56, 56, 56
        2496 => x"38383939",		-- colors: 56, 56, 57, 57
        2497 => x"39393939",		-- colors: 57, 57, 57, 57
        2498 => x"38383838",		-- colors: 56, 56, 56, 56
        2499 => x"38383838",		-- colors: 56, 56, 56, 56
        2500 => x"38393939",		-- colors: 56, 57, 57, 57
        2501 => x"39393939",		-- colors: 57, 57, 57, 57
        2502 => x"39383838",		-- colors: 57, 56, 56, 56
        2503 => x"38393938",		-- colors: 56, 57, 57, 56
        2504 => x"38393A39",		-- colors: 56, 57, 58, 57
        2505 => x"3A3A3A3A",		-- colors: 58, 58, 58, 58
        2506 => x"38383838",		-- colors: 56, 56, 56, 56
        2507 => x"38383839",		-- colors: 56, 56, 56, 57
        2508 => x"3939393A",		-- colors: 57, 57, 57, 58
        2509 => x"3A3A393A",		-- colors: 58, 58, 57, 58
        2510 => x"3A383838",		-- colors: 58, 56, 56, 56
        2511 => x"38393939",		-- colors: 56, 57, 57, 57
        2512 => x"39393A3A",		-- colors: 57, 57, 58, 58
        2513 => x"3A3A3A3A",		-- colors: 58, 58, 58, 58
        2514 => x"38383838",		-- colors: 56, 56, 56, 56
        2515 => x"38383939",		-- colors: 56, 56, 57, 57
        2516 => x"3938393A",		-- colors: 57, 56, 57, 58
        2517 => x"3A3A3A38",		-- colors: 58, 58, 58, 56
        2518 => x"38383838",		-- colors: 56, 56, 56, 56
        2519 => x"38393938",		-- colors: 56, 57, 57, 56
        2520 => x"383B3B3A",		-- colors: 56, 59, 59, 58
        2521 => x"3A383838",		-- colors: 58, 56, 56, 56
        2522 => x"38383838",		-- colors: 56, 56, 56, 56
        2523 => x"38383838",		-- colors: 56, 56, 56, 56
        2524 => x"3B3B3B3B",		-- colors: 59, 59, 59, 59
        2525 => x"3B383838",		-- colors: 59, 56, 56, 56
        2526 => x"38383838",		-- colors: 56, 56, 56, 56
        2527 => x"38383838",		-- colors: 56, 56, 56, 56
        2528 => x"3A3B3B3B",		-- colors: 58, 59, 59, 59
        2529 => x"3B3B383A",		-- colors: 59, 59, 56, 58
        2530 => x"38383838",		-- colors: 56, 56, 56, 56
        2531 => x"3838383A",		-- colors: 56, 56, 56, 58
        2532 => x"3A3A3B3B",		-- colors: 58, 58, 59, 59
        2533 => x"3B3B3A3A",		-- colors: 59, 59, 58, 58
        2534 => x"3A383838",		-- colors: 58, 56, 56, 56
        2535 => x"38383A3A",		-- colors: 56, 56, 58, 58
        2536 => x"3B3B3A3A",		-- colors: 59, 59, 58, 58
        2537 => x"3A3B3A3A",		-- colors: 58, 59, 58, 58
        2538 => x"38383838",		-- colors: 56, 56, 56, 56
        2539 => x"38383B3B",		-- colors: 56, 56, 59, 59
        2540 => x"3B3B3B3B",		-- colors: 59, 59, 59, 59
        2541 => x"3B3B3B38",		-- colors: 59, 59, 59, 56
        2542 => x"38383838",		-- colors: 56, 56, 56, 56
        2543 => x"39383B3B",		-- colors: 57, 56, 59, 59
        2544 => x"3B3B3B3B",		-- colors: 59, 59, 59, 59
        2545 => x"3B3B3B38",		-- colors: 59, 59, 59, 56
        2546 => x"38383838",		-- colors: 56, 56, 56, 56
        2547 => x"39393A3A",		-- colors: 57, 57, 58, 58
        2548 => x"3A3A3A3A",		-- colors: 58, 58, 58, 58
        2549 => x"3A3A3A3A",		-- colors: 58, 58, 58, 58
        2550 => x"38383838",		-- colors: 56, 56, 56, 56
        2551 => x"39383838",		-- colors: 57, 56, 56, 56
        2552 => x"38383838",		-- colors: 56, 56, 56, 56
        2553 => x"39393838",		-- colors: 57, 57, 56, 56
        2554 => x"38383838",		-- colors: 56, 56, 56, 56
        2555 => x"38383838",		-- colors: 56, 56, 56, 56
        2556 => x"38383838",		-- colors: 56, 56, 56, 56
        2557 => x"39393938",		-- colors: 57, 57, 57, 56
        2558 => x"38383838",		-- colors: 56, 56, 56, 56
		  --heart
		  --  sprite 0
        2559 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
        2560 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
        2561 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
        2562 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
        2563 => x"3C3C3D3D",		-- colors: 60, 60, 61, 61
        2564 => x"3D3D3D3D",		-- colors: 61, 61, 61, 61
        2565 => x"3C3D3D3D",		-- colors: 60, 61, 61, 61
        2566 => x"3D3D3D3C",		-- colors: 61, 61, 61, 60
        2567 => x"3C3D3D3E",		-- colors: 60, 61, 61, 62
        2568 => x"3E3E3E3D",		-- colors: 62, 62, 62, 61
        2569 => x"3D3D3E3E",		-- colors: 61, 61, 62, 62
        2570 => x"3E3E3D3D",		-- colors: 62, 62, 61, 61
        2571 => x"3D3D3E3E",		-- colors: 61, 61, 62, 62
        2572 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
        2573 => x"3D3E3E3E",		-- colors: 61, 62, 62, 62
        2574 => x"3E3E3E3D",		-- colors: 62, 62, 62, 61
        2575 => x"3D3E3E3E",		-- colors: 61, 62, 62, 62
        2576 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
        2577 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
        2578 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
        2579 => x"3D3E3E3E",		-- colors: 61, 62, 62, 62
        2580 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
        2581 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
        2582 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
        2583 => x"3D3E3E3E",		-- colors: 61, 62, 62, 62
        2584 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
        2585 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
        2586 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
        2587 => x"3D3E3E3E",		-- colors: 61, 62, 62, 62
        2588 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
        2589 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
        2590 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
        2591 => x"3D3D3E3E",		-- colors: 61, 61, 62, 62
        2592 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
        2593 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
        2594 => x"3E3E3E3D",		-- colors: 62, 62, 62, 61
        2595 => x"3C3D3E3E",		-- colors: 60, 61, 62, 62
        2596 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
        2597 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
        2598 => x"3E3E3E3D",		-- colors: 62, 62, 62, 61
        2599 => x"3C3D3D3E",		-- colors: 60, 61, 61, 62
        2600 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
        2601 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
        2602 => x"3E3E3D3D",		-- colors: 62, 62, 61, 61
        2603 => x"3C3C3D3D",		-- colors: 60, 60, 61, 61
        2604 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
        2605 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
        2606 => x"3E3D3D3C",		-- colors: 62, 61, 61, 60
        2607 => x"3C3C3C3D",		-- colors: 60, 60, 60, 61
        2608 => x"3D3D3E3E",		-- colors: 61, 61, 62, 62
        2609 => x"3E3E3E3D",		-- colors: 62, 62, 62, 61
        2610 => x"3D3D3C3C",		-- colors: 61, 61, 60, 60
        2611 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
        2612 => x"3C3D3D3E",		-- colors: 60, 61, 61, 62
        2613 => x"3E3E3D3D",		-- colors: 62, 62, 61, 61
        2614 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
        2615 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
        2616 => x"3C3C3D3D",		-- colors: 60, 60, 61, 61
        2617 => x"3E3D3D3C",		-- colors: 62, 61, 61, 60
        2618 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
        2619 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
        2620 => x"3C3C3C3D",		-- colors: 60, 60, 60, 61
        2621 => x"3D3D3C3C",		-- colors: 61, 61, 60, 60
        2622 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60

				-----------------------------------------------
		--****  MAP  ****
        6992 => x"00000016", -- pedding
        6993 => x"00000016", -- pedding
        6994 => x"00000016", -- pedding
        6995 => x"00000016", -- pedding
        6996 => x"00000016", -- pedding
        6997 => x"00000016", -- pedding
        6998 => x"00000016", -- pedding
        6999 => x"00000016", -- pedding
        7000 => x"00000016", -- pedding
        7001 => x"00000016", -- pedding
        7002 => x"00000016", -- pedding
        7003 => x"00000016", -- pedding
        7004 => x"00000016", -- pedding
        7005 => x"00000016", -- pedding
        7006 => x"00000016", -- pedding
        7007 => x"00000016", -- pedding
        7008 => x"00000016", -- pedding
        7009 => x"00000016", -- pedding
        7010 => x"00000016", -- pedding
        7011 => x"00000016", -- pedding
        7012 => x"00000016", -- pedding
        7013 => x"00000016", -- pedding
        7014 => x"00000016", -- pedding
        7015 => x"00000016", -- pedding
        7016 => x"00000016", -- pedding
        7017 => x"00000016", -- pedding
        7018 => x"00000016", -- pedding
        7019 => x"00000016", -- pedding
        7020 => x"00000016", -- pedding
        7021 => x"00000016", -- pedding
        7022 => x"00000016", -- pedding
        7023 => x"00000016", -- pedding
        7024 => x"00000016", -- pedding
        7025 => x"00000016", -- pedding
        7026 => x"00000016", -- pedding
        7027 => x"00000016", -- pedding
        7028 => x"00000016", -- pedding
        7029 => x"00000016", -- pedding
        7030 => x"00000016", -- pedding
        7031 => x"00000016", -- pedding
        7032 => x"00000016", -- pedding
        7033 => x"00000016", -- pedding
        7034 => x"00000016", -- pedding
        7035 => x"00000016", -- pedding
        7036 => x"00000016", -- pedding
        7037 => x"00000016", -- pedding
        7038 => x"00000016", -- pedding
        7039 => x"00000016", -- pedding
        7040 => x"00000016", -- pedding
        7041 => x"00000016", -- pedding
        7042 => x"00000016", -- pedding
        7043 => x"00000016", -- pedding
        7044 => x"00000016", -- pedding
        7045 => x"00000016", -- pedding
        7046 => x"00000016", -- pedding
        7047 => x"00000016", -- pedding
        7048 => x"00000016", -- pedding
        7049 => x"00000016", -- pedding
        7050 => x"00000016", -- pedding
        7051 => x"00000016", -- pedding
        7052 => x"00000016", -- pedding
        7053 => x"00000016", -- pedding
        7054 => x"00000016", -- pedding
        7055 => x"00000016", -- pedding
        7056 => x"00000016", -- pedding
        7057 => x"00000016", -- pedding
        7058 => x"00000016", -- pedding
        7059 => x"00000016", -- pedding
        7060 => x"00000016", -- pedding
        7061 => x"00000016", -- pedding
        7062 => x"00000016", -- pedding
        7063 => x"00000016", -- pedding
        7064 => x"00000016", -- pedding
        7065 => x"00000016", -- pedding
        7066 => x"00000016", -- pedding
        7067 => x"00000016", -- pedding
        7068 => x"00000016", -- pedding
        7069 => x"00000016", -- pedding
        7070 => x"00000016", -- pedding
        7071 => x"00000016", -- pedding
        7072 => x"00000016", -- pedding
        7073 => x"00000016", -- pedding
        7074 => x"00000016", -- pedding
        7075 => x"00000016", -- pedding
        7076 => x"00000016", -- pedding
        7077 => x"00000016", -- pedding
        7078 => x"00000016", -- pedding
        7079 => x"00000016", -- pedding
        7080 => x"00000016", -- pedding
        7081 => x"00000016", -- pedding
        7082 => x"00000016", -- pedding
        7083 => x"00000016", -- pedding
        7084 => x"00000016", -- pedding
        7085 => x"00000016", -- pedding
        7086 => x"00000016", -- pedding
        7087 => x"00000016", -- pedding
        7088 => x"00000016", -- pedding
        7089 => x"00000016", -- pedding
        7090 => x"00000016", -- pedding
        7091 => x"00000016", -- pedding
        7092 => x"00000016", -- pedding
        7093 => x"00000016", -- pedding
        7094 => x"00000016", -- pedding
        7095 => x"00000016", -- pedding
        7096 => x"00000016", -- pedding
        7097 => x"00000016", -- pedding
        7098 => x"00000016", -- pedding
        7099 => x"00000016", -- pedding
        7100 => x"00000016", -- pedding
        7101 => x"00000016", -- pedding
        7102 => x"00000016", -- pedding
        7103 => x"00000016", -- pedding
        7104 => x"00000016", -- pedding
        7105 => x"00000016", -- pedding
        7106 => x"00000016", -- pedding
        7107 => x"00000016", -- pedding
        7108 => x"00000016", -- pedding
        7109 => x"00000016", -- pedding
        7110 => x"00000016", -- pedding
        7111 => x"00000016", -- pedding
        7112 => x"00000016", -- pedding
        7113 => x"00000016", -- pedding
        7114 => x"00000016", -- pedding
        7115 => x"00000016", -- pedding
        7116 => x"00000016", -- pedding
        7117 => x"00000016", -- pedding
        7118 => x"00000016", -- pedding
        7119 => x"00000016", -- pedding
        7120 => x"00000016", -- pedding
        7121 => x"00000016", -- pedding
        7122 => x"00000016", -- pedding
        7123 => x"00000016", -- pedding
        7124 => x"00000016", -- header
        7125 => x"00000016", -- header
        7126 => x"00000016", -- header
        7127 => x"00000016", -- header
        7128 => x"00000016", -- header
        7129 => x"00000016", -- header
        7130 => x"00000016", -- header
        7131 => x"00000016", -- header
        7132 => x"00000016", -- header
        7133 => x"00000016", -- header
        7134 => x"00000016", -- header
        7135 => x"00000016", -- header
        7136 => x"00000016", -- header
        7137 => x"00000016", -- header
        7138 => x"00000016", -- header
        7139 => x"00000016", -- header
        7140 => x"00000016", -- pedding
        7141 => x"00000016", -- pedding
        7142 => x"00000016", -- pedding
        7143 => x"00000016", -- pedding
        7144 => x"00000016", -- pedding
        7145 => x"00000016", -- pedding
        7146 => x"00000016", -- pedding
        7147 => x"00000016", -- pedding
        7148 => x"00000016", -- pedding
        7149 => x"00000016", -- pedding
        7150 => x"00000016", -- pedding
        7151 => x"00000016", -- pedding
        7152 => x"00000016", -- pedding
        7153 => x"00000016", -- pedding
        7154 => x"00000016", -- pedding
        7155 => x"00000016", -- pedding
        7156 => x"00000016", -- pedding
        7157 => x"00000016", -- pedding
        7158 => x"00000016", -- pedding
        7159 => x"00000016", -- pedding
        7160 => x"00000016", -- pedding
        7161 => x"00000016", -- pedding
        7162 => x"00000016", -- pedding
        7163 => x"00000016", -- pedding
        7164 => x"00000016", -- header
        7165 => x"00000016", -- header
        7166 => x"00000016", -- header
        7167 => x"00000016", -- header
        7168 => x"00000016", -- header
        7169 => x"00000016", -- header
        7170 => x"00000016", -- header
        7171 => x"00000016", -- header
        7172 => x"00000016", -- header
        7173 => x"00000016", -- header
        7174 => x"00000016", -- header
        7175 => x"00000016", -- header
        7176 => x"00000016", -- header
        7177 => x"00000016", -- header
        7178 => x"00000016", -- header
        7179 => x"00000016", -- header
        7180 => x"00000016", -- pedding
        7181 => x"00000016", -- pedding
        7182 => x"00000016", -- pedding
        7183 => x"00000016", -- pedding
        7184 => x"00000016", -- pedding
        7185 => x"00000016", -- pedding
        7186 => x"00000016", -- pedding
        7187 => x"00000016", -- pedding
        7188 => x"00000016", -- pedding
        7189 => x"00000016", -- pedding
        7190 => x"00000016", -- pedding
        7191 => x"00000016", -- pedding
        7192 => x"00000016", -- pedding
        7193 => x"00000016", -- pedding
        7194 => x"00000016", -- pedding
        7195 => x"00000016", -- pedding
        7196 => x"00000016", -- pedding
        7197 => x"00000016", -- pedding
        7198 => x"00000016", -- pedding
        7199 => x"00000016", -- pedding
        7200 => x"00000016", -- pedding
        7201 => x"00000016", -- pedding
        7202 => x"00000016", -- pedding
        7203 => x"00000016", -- pedding
        7204 => x"00000016", -- header
        7205 => x"00000016", -- header
        7206 => x"00000016", -- header
        7207 => x"00000016", -- header
        7208 => x"00000016", -- header
        7209 => x"00000016", -- header
        7210 => x"00000016", -- header
        7211 => x"00000016", -- header
        7212 => x"00000016", -- header
        7213 => x"00000016", -- header
        7214 => x"00000016", -- header
        7215 => x"00000016", -- header
        7216 => x"00000016", -- header
        7217 => x"00000016", -- header
        7218 => x"00000016", -- header
        7219 => x"00000016", -- header
        7220 => x"00000016", -- pedding
        7221 => x"00000016", -- pedding
        7222 => x"00000016", -- pedding
        7223 => x"00000016", -- pedding
        7224 => x"00000016", -- pedding
        7225 => x"00000016", -- pedding
        7226 => x"00000016", -- pedding
        7227 => x"00000016", -- pedding
        7228 => x"00000016", -- pedding
        7229 => x"00000016", -- pedding
        7230 => x"00000016", -- pedding
        7231 => x"00000016", -- pedding
        7232 => x"00000016", -- pedding
        7233 => x"00000016", -- pedding
        7234 => x"00000016", -- pedding
        7235 => x"00000016", -- pedding
        7236 => x"00000016", -- pedding
        7237 => x"00000016", -- pedding
        7238 => x"00000016", -- pedding
        7239 => x"00000016", -- pedding
        7240 => x"00000016", -- pedding
        7241 => x"00000016", -- pedding
        7242 => x"00000016", -- pedding
        7243 => x"00000016", -- pedding
        7244 => x"00000016", -- header
        7245 => x"00000016", -- header
        7246 => x"00000016", -- header
        7247 => x"00000016", -- header
        7248 => x"00000016", -- header
        7249 => x"00000016", -- header
        7250 => x"00000016", -- header
        7251 => x"00000016", -- header
        7252 => x"00000016", -- header
        7253 => x"00000016", -- header
        7254 => x"00000016", -- header
        7255 => x"00000016", -- header
        7256 => x"00000016", -- header
        7257 => x"00000016", -- header
        7258 => x"00000016", -- header
        7259 => x"00000016", -- header
        7260 => x"00000016", -- pedding
        7261 => x"00000016", -- pedding
        7262 => x"00000016", -- pedding
        7263 => x"00000016", -- pedding
        7264 => x"00000016", -- pedding
        7265 => x"00000016", -- pedding
        7266 => x"00000016", -- pedding
        7267 => x"00000016", -- pedding
        7268 => x"00000016", -- pedding
        7269 => x"00000016", -- pedding
        7270 => x"00000016", -- pedding
        7271 => x"00000016", -- pedding
        7272 => x"00000016", -- pedding
        7273 => x"00000016", -- pedding
        7274 => x"00000016", -- pedding
        7275 => x"00000016", -- pedding
        7276 => x"00000016", -- pedding
        7277 => x"00000016", -- pedding
        7278 => x"00000016", -- pedding
        7279 => x"00000016", -- pedding
        7280 => x"00000016", -- pedding
        7281 => x"00000016", -- pedding
        7282 => x"00000016", -- pedding
        7283 => x"00000016", -- pedding
        7284 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7285 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7286 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7287 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7288 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7289 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7290 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7291 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7292 => x"00000001", -- z: 0 rot: 0 ptr: 319
        7293 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7294 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7295 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7296 => x"00000001", -- z: 0 rot: 0 ptr: 319
        7297 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7298 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7299 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7300 => x"00000016", -- pedding
        7301 => x"00000016", -- pedding
        7302 => x"00000016", -- pedding
        7303 => x"00000016", -- pedding
        7304 => x"00000016", -- pedding
        7305 => x"00000016", -- pedding
        7306 => x"00000016", -- pedding
        7307 => x"00000016", -- pedding
        7308 => x"00000016", -- pedding
        7309 => x"00000016", -- pedding
        7310 => x"00000016", -- pedding
        7311 => x"00000016", -- pedding
        7312 => x"00000016", -- pedding
        7313 => x"00000016", -- pedding
        7314 => x"00000016", -- pedding
        7315 => x"00000016", -- pedding
        7316 => x"00000016", -- pedding
        7317 => x"00000016", -- pedding
        7318 => x"00000016", -- pedding
        7319 => x"00000016", -- pedding
        7320 => x"00000016", -- pedding
        7321 => x"00000016", -- pedding
        7322 => x"00000016", -- pedding
        7323 => x"00000016", -- pedding
        7324 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7325 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7326 => x"00000003", -- z: 0 rot: 0 ptr: 447
        7327 => x"00000005", -- z: 0 rot: 0 ptr: 575
        7328 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7329 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7330 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7331 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7332 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7333 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7334 => x"00000001", -- z: 0 rot: 0 ptr: 319
        7335 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7336 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7337 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7338 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7339 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7340 => x"00000016", -- pedding
        7341 => x"00000016", -- pedding
        7342 => x"00000016", -- pedding
        7343 => x"00000016", -- pedding
        7344 => x"00000016", -- pedding
        7345 => x"00000016", -- pedding
        7346 => x"00000016", -- pedding
        7347 => x"00000016", -- pedding
        7348 => x"00000016", -- pedding
        7349 => x"00000016", -- pedding
        7350 => x"00000016", -- pedding
        7351 => x"00000016", -- pedding
        7352 => x"00000016", -- pedding
        7353 => x"00000016", -- pedding
        7354 => x"00000016", -- pedding
        7355 => x"00000016", -- pedding
        7356 => x"00000016", -- pedding
        7357 => x"00000016", -- pedding
        7358 => x"00000016", -- pedding
        7359 => x"00000016", -- pedding
        7360 => x"00000016", -- pedding
        7361 => x"00000016", -- pedding
        7362 => x"00000016", -- pedding
        7363 => x"00000016", -- pedding
        7364 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7365 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7366 => x"00000015", -- z: 0 rot: 0 ptr: 831
        7367 => x"00000017", -- z: 0 rot: 0 ptr: 959
        7368 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7369 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7370 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7371 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7372 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7373 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7374 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7375 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7376 => x"00000001", -- z: 0 rot: 0 ptr: 319
        7377 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7378 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7379 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7380 => x"00000016", -- pedding
        7381 => x"00000016", -- pedding
        7382 => x"00000016", -- pedding
        7383 => x"00000016", -- pedding
        7384 => x"00000016", -- pedding
        7385 => x"00000016", -- pedding
        7386 => x"00000016", -- pedding
        7387 => x"00000016", -- pedding
        7388 => x"00000016", -- pedding
        7389 => x"00000016", -- pedding
        7390 => x"00000016", -- pedding
        7391 => x"00000016", -- pedding
        7392 => x"00000016", -- pedding
        7393 => x"00000016", -- pedding
        7394 => x"00000016", -- pedding
        7395 => x"00000016", -- pedding
        7396 => x"00000016", -- pedding
        7397 => x"00000016", -- pedding
        7398 => x"00000016", -- pedding
        7399 => x"00000016", -- pedding
        7400 => x"00000016", -- pedding
        7401 => x"00000016", -- pedding
        7402 => x"00000016", -- pedding
        7403 => x"00000016", -- pedding
        7404 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7405 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7406 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7407 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7408 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7409 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7410 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7411 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7412 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7413 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7414 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7415 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7416 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7417 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7418 => x"00000024", -- z: 0 rot: 0 ptr: 1023
        7419 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7420 => x"00000016", -- pedding
        7421 => x"00000016", -- pedding
        7422 => x"00000016", -- pedding
        7423 => x"00000016", -- pedding
        7424 => x"00000016", -- pedding
        7425 => x"00000016", -- pedding
        7426 => x"00000016", -- pedding
        7427 => x"00000016", -- pedding
        7428 => x"00000016", -- pedding
        7429 => x"00000016", -- pedding
        7430 => x"00000016", -- pedding
        7431 => x"00000016", -- pedding
        7432 => x"00000016", -- pedding
        7433 => x"00000016", -- pedding
        7434 => x"00000016", -- pedding
        7435 => x"00000016", -- pedding
        7436 => x"00000016", -- pedding
        7437 => x"00000016", -- pedding
        7438 => x"00000016", -- pedding
        7439 => x"00000016", -- pedding
        7440 => x"00000016", -- pedding
        7441 => x"00000016", -- pedding
        7442 => x"00000016", -- pedding
        7443 => x"00000016", -- pedding
        7444 => x"00000025", -- z: 0 rot: 0 ptr: 1087
        7445 => x"00000025", -- z: 0 rot: 0 ptr: 1087
        7446 => x"00000025", -- z: 0 rot: 0 ptr: 1087
        7447 => x"00000025", -- z: 0 rot: 0 ptr: 1087
        7448 => x"00000025", -- z: 0 rot: 0 ptr: 1087
        7449 => x"00000025", -- z: 0 rot: 0 ptr: 1087
        7450 => x"00000025", -- z: 0 rot: 0 ptr: 1087
        7451 => x"00000025", -- z: 0 rot: 0 ptr: 1087
        7452 => x"00000025", -- z: 0 rot: 0 ptr: 1087
        7453 => x"00000025", -- z: 0 rot: 0 ptr: 1087
        7454 => x"00000025", -- z: 0 rot: 0 ptr: 1087
        7455 => x"00000025", -- z: 0 rot: 0 ptr: 1087
        7456 => x"00000025", -- z: 0 rot: 0 ptr: 1087
        7457 => x"00000025", -- z: 0 rot: 0 ptr: 1087
        7458 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7459 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7460 => x"00000016", -- pedding
        7461 => x"00000016", -- pedding
        7462 => x"00000016", -- pedding
        7463 => x"00000016", -- pedding
        7464 => x"00000016", -- pedding
        7465 => x"00000016", -- pedding
        7466 => x"00000016", -- pedding
        7467 => x"00000016", -- pedding
        7468 => x"00000016", -- pedding
        7469 => x"00000016", -- pedding
        7470 => x"00000016", -- pedding
        7471 => x"00000016", -- pedding
        7472 => x"00000016", -- pedding
        7473 => x"00000016", -- pedding
        7474 => x"00000016", -- pedding
        7475 => x"00000016", -- pedding
        7476 => x"00000016", -- pedding
        7477 => x"00000016", -- pedding
        7478 => x"00000016", -- pedding
        7479 => x"00000016", -- pedding
        7480 => x"00000016", -- pedding
        7481 => x"00000016", -- pedding
        7482 => x"00000016", -- pedding
        7483 => x"00000016", -- pedding
        7484 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7485 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7486 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7487 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7488 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7489 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7490 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7491 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7492 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7493 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7494 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7495 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7496 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7497 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7498 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7499 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7500 => x"00000016", -- pedding
        7501 => x"00000016", -- pedding
        7502 => x"00000016", -- pedding
        7503 => x"00000016", -- pedding
        7504 => x"00000016", -- pedding
        7505 => x"00000016", -- pedding
        7506 => x"00000016", -- pedding
        7507 => x"00000016", -- pedding
        7508 => x"00000016", -- pedding
        7509 => x"00000016", -- pedding
        7510 => x"00000016", -- pedding
        7511 => x"00000016", -- pedding
        7512 => x"00000016", -- pedding
        7513 => x"00000016", -- pedding
        7514 => x"00000016", -- pedding
        7515 => x"00000016", -- pedding
        7516 => x"00000016", -- pedding
        7517 => x"00000016", -- pedding
        7518 => x"00000016", -- pedding
        7519 => x"00000016", -- pedding
        7520 => x"00000016", -- pedding
        7521 => x"00000016", -- pedding
        7522 => x"00000016", -- pedding
        7523 => x"00000016", -- pedding
        7524 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7525 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7526 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7527 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7528 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7529 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7530 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7531 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7532 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7533 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7534 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7535 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7536 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7537 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7538 => x"00000013", -- z: 0 rot: 0 ptr: 703
        7539 => x"00000013", -- z: 0 rot: 0 ptr: 703
        7540 => x"00000016", -- pedding
        7541 => x"00000016", -- pedding
        7542 => x"00000016", -- pedding
        7543 => x"00000016", -- pedding
        7544 => x"00000016", -- pedding
        7545 => x"00000016", -- pedding
        7546 => x"00000016", -- pedding
        7547 => x"00000016", -- pedding
        7548 => x"00000016", -- pedding
        7549 => x"00000016", -- pedding
        7550 => x"00000016", -- pedding
        7551 => x"00000016", -- pedding
        7552 => x"00000016", -- pedding
        7553 => x"00000016", -- pedding
        7554 => x"00000016", -- pedding
        7555 => x"00000016", -- pedding
        7556 => x"00000016", -- pedding
        7557 => x"00000016", -- pedding
        7558 => x"00000016", -- pedding
        7559 => x"00000016", -- pedding
        7560 => x"00000016", -- pedding
        7561 => x"00000016", -- pedding
        7562 => x"00000016", -- pedding
        7563 => x"00000016", -- pedding
        7564 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7565 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7566 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7567 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7568 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7569 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7570 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7571 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7572 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7573 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7574 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7575 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7576 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7577 => x"00000037", -- z: 0 rot: 0 ptr: 1471
        7578 => x"00000013", -- z: 0 rot: 0 ptr: 703
        7579 => x"00000013", -- z: 0 rot: 0 ptr: 703
        7580 => x"00000016", -- pedding
        7581 => x"00000016", -- pedding
        7582 => x"00000016", -- pedding
        7583 => x"00000016", -- pedding
        7584 => x"00000016", -- pedding
        7585 => x"00000016", -- pedding
        7586 => x"00000016", -- pedding
        7587 => x"00000016", -- pedding
        7588 => x"00000016", -- pedding
        7589 => x"00000016", -- pedding
        7590 => x"00000016", -- pedding
        7591 => x"00000016", -- pedding
        7592 => x"00000016", -- pedding
        7593 => x"00000016", -- pedding
        7594 => x"00000016", -- pedding
        7595 => x"00000016", -- pedding
        7596 => x"00000016", -- pedding
        7597 => x"00000016", -- pedding
        7598 => x"00000016", -- pedding
        7599 => x"00000016", -- pedding
        7600 => x"00000016", -- pedding
        7601 => x"00000016", -- pedding
        7602 => x"00000016", -- pedding
        7603 => x"00000016", -- pedding
        7604 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7605 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7606 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7607 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7608 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7609 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7610 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7611 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7612 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7613 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7614 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7615 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7616 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7617 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7618 => x"00000013", -- z: 0 rot: 0 ptr: 703
        7619 => x"00000013", -- z: 0 rot: 0 ptr: 703
        7620 => x"00000016", -- pedding
        7621 => x"00000016", -- pedding
        7622 => x"00000016", -- pedding
        7623 => x"00000016", -- pedding
        7624 => x"00000016", -- pedding
        7625 => x"00000016", -- pedding
        7626 => x"00000016", -- pedding
        7627 => x"00000016", -- pedding
        7628 => x"00000016", -- pedding
        7629 => x"00000016", -- pedding
        7630 => x"00000016", -- pedding
        7631 => x"00000016", -- pedding
        7632 => x"00000016", -- pedding
        7633 => x"00000016", -- pedding
        7634 => x"00000016", -- pedding
        7635 => x"00000016", -- pedding
        7636 => x"00000016", -- pedding
        7637 => x"00000016", -- pedding
        7638 => x"00000016", -- pedding
        7639 => x"00000016", -- pedding
        7640 => x"00000016", -- pedding
        7641 => x"00000016", -- pedding
        7642 => x"00000016", -- pedding
        7643 => x"00000016", -- pedding
        7644 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7645 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7646 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7647 => x"00000092", -- z: 0 rot: 0 ptr: 3455
        7648 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7649 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7650 => x"00000092", -- z: 0 rot: 0 ptr: 3455
        7651 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7652 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7653 => x"00000092", -- z: 0 rot: 0 ptr: 3455
        7654 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7655 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7656 => x"00000092", -- z: 0 rot: 0 ptr: 3455
        7657 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7658 => x"00000013", -- z: 0 rot: 0 ptr: 703
        7659 => x"00000013", -- z: 0 rot: 0 ptr: 703
        7660 => x"00000016", -- pedding
        7661 => x"00000016", -- pedding
        7662 => x"00000016", -- pedding
        7663 => x"00000016", -- pedding
        7664 => x"00000016", -- pedding
        7665 => x"00000016", -- pedding
        7666 => x"00000016", -- pedding
        7667 => x"00000016", -- pedding
        7668 => x"00000016", -- pedding
        7669 => x"00000016", -- pedding
        7670 => x"00000016", -- pedding
        7671 => x"00000016", -- pedding
        7672 => x"00000016", -- pedding
        7673 => x"00000016", -- pedding
        7674 => x"00000016", -- pedding
        7675 => x"00000016", -- pedding
        7676 => x"00000016", -- pedding
        7677 => x"00000016", -- pedding
        7678 => x"00000016", -- pedding
        7679 => x"00000016", -- pedding
        7680 => x"00000016", -- pedding
        7681 => x"00000016", -- pedding
        7682 => x"00000016", -- pedding
        7683 => x"00000016", -- pedding
        7684 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7685 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7686 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7687 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7688 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7689 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7690 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7691 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7692 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7693 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7694 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7695 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7696 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7697 => x"00000002", -- z: 0 rot: 0 ptr: 383
        7698 => x"00000013", -- z: 0 rot: 0 ptr: 703
        7699 => x"00000013", -- z: 0 rot: 0 ptr: 703
        7700 => x"00000016", -- pedding
        7701 => x"00000016", -- pedding
        7702 => x"00000016", -- pedding
        7703 => x"00000016", -- pedding
        7704 => x"00000016", -- pedding
        7705 => x"00000016", -- pedding
        7706 => x"00000016", -- pedding
        7707 => x"00000016", -- pedding
        7708 => x"00000016", -- pedding
        7709 => x"00000016", -- pedding
        7710 => x"00000016", -- pedding
        7711 => x"00000016", -- pedding
        7712 => x"00000016", -- pedding
        7713 => x"00000016", -- pedding
        7714 => x"00000016", -- pedding
        7715 => x"00000016", -- pedding
        7716 => x"00000016", -- pedding
        7717 => x"00000016", -- pedding
        7718 => x"00000016", -- pedding
        7719 => x"00000016", -- pedding
        7720 => x"00000016", -- pedding
        7721 => x"00000016", -- pedding
        7722 => x"00000016", -- pedding
        7723 => x"00000016", -- pedding
        7724 => x"00000016", -- pedding
        7725 => x"00000016", -- pedding
        7726 => x"00000016", -- pedding
        7727 => x"00000016", -- pedding
        7728 => x"00000016", -- pedding
        7729 => x"00000016", -- pedding
        7730 => x"00000016", -- pedding
        7731 => x"00000016", -- pedding
        7732 => x"00000016", -- pedding
        7733 => x"00000016", -- pedding
        7734 => x"00000016", -- pedding
        7735 => x"00000016", -- pedding
        7736 => x"00000016", -- pedding
        7737 => x"00000016", -- pedding
        7738 => x"00000016", -- pedding
        7739 => x"00000016", -- pedding
        7740 => x"00000016", -- pedding
        7741 => x"00000016", -- pedding
        7742 => x"00000016", -- pedding
        7743 => x"00000016", -- pedding
        7744 => x"00000016", -- pedding
        7745 => x"00000016", -- pedding
        7746 => x"00000016", -- pedding
        7747 => x"00000016", -- pedding
        7748 => x"00000016", -- pedding
        7749 => x"00000016", -- pedding
        7750 => x"00000016", -- pedding
        7751 => x"00000016", -- pedding
        7752 => x"00000016", -- pedding
        7753 => x"00000016", -- pedding
        7754 => x"00000016", -- pedding
        7755 => x"00000016", -- pedding
        7756 => x"00000016", -- pedding
        7757 => x"00000016", -- pedding
        7758 => x"00000016", -- pedding
        7759 => x"00000016", -- pedding
        7760 => x"00000016", -- pedding
        7761 => x"00000016", -- pedding
        7762 => x"00000016", -- pedding
        7763 => x"00000016", -- pedding
        7764 => x"00000016", -- pedding
        7765 => x"00000016", -- pedding
        7766 => x"00000016", -- pedding
        7767 => x"00000016", -- pedding
        7768 => x"00000016", -- pedding
        7769 => x"00000016", -- pedding
        7770 => x"00000016", -- pedding
        7771 => x"00000016", -- pedding
        7772 => x"00000016", -- pedding
        7773 => x"00000016", -- pedding
        7774 => x"00000016", -- pedding
        7775 => x"00000016", -- pedding
        7776 => x"00000016", -- pedding
        7777 => x"00000016", -- pedding
        7778 => x"00000016", -- pedding
        7779 => x"00000016", -- pedding
        7780 => x"00000016", -- pedding
        7781 => x"00000016", -- pedding
        7782 => x"00000016", -- pedding
        7783 => x"00000016", -- pedding
        7784 => x"00000016", -- pedding
        7785 => x"00000016", -- pedding
        7786 => x"00000016", -- pedding
        7787 => x"00000016", -- pedding
        7788 => x"00000016", -- pedding
        7789 => x"00000016", -- pedding
        7790 => x"00000016", -- pedding
        7791 => x"00000016", -- pedding
        7792 => x"00000016", -- pedding
        7793 => x"00000016", -- pedding
        7794 => x"00000016", -- pedding
        7795 => x"00000016", -- pedding
        7796 => x"00000016", -- pedding
        7797 => x"00000016", -- pedding
        7798 => x"00000016", -- pedding
        7799 => x"00000016", -- pedding
        7800 => x"00000016", -- pedding
        7801 => x"00000016", -- pedding
        7802 => x"00000016", -- pedding
        7803 => x"00000016", -- pedding
        7804 => x"00000016", -- pedding
        7805 => x"00000016", -- pedding
        7806 => x"00000016", -- pedding
        7807 => x"00000016", -- pedding
        7808 => x"00000016", -- pedding
        7809 => x"00000016", -- pedding
        7810 => x"00000016", -- pedding
        7811 => x"00000016", -- pedding
        7812 => x"00000016", -- pedding
        7813 => x"00000016", -- pedding
        7814 => x"00000016", -- pedding
        7815 => x"00000016", -- pedding
        7816 => x"00000016", -- pedding
        7817 => x"00000016", -- pedding
        7818 => x"00000016", -- pedding
        7819 => x"00000016", -- pedding
        7820 => x"00000016", -- pedding
        7821 => x"00000016", -- pedding
        7822 => x"00000016", -- pedding
        7823 => x"00000016", -- pedding
        7824 => x"00000016", -- pedding
        7825 => x"00000016", -- pedding
        7826 => x"00000016", -- pedding
        7827 => x"00000016", -- pedding
        7828 => x"00000016", -- pedding
        7829 => x"00000016", -- pedding
        7830 => x"00000016", -- pedding
        7831 => x"00000016", -- pedding
        7832 => x"00000016", -- pedding
        7833 => x"00000016", -- pedding
        7834 => x"00000016", -- pedding
        7835 => x"00000016", -- pedding
        7836 => x"00000016", -- pedding
        7837 => x"00000016", -- pedding
        7838 => x"00000016", -- pedding
        7839 => x"00000016", -- pedding
        7840 => x"00000016", -- pedding
        7841 => x"00000016", -- pedding
        7842 => x"00000016", -- pedding
        7843 => x"00000016", -- pedding
        7844 => x"00000016", -- pedding
        7845 => x"00000016", -- pedding
        7846 => x"00000016", -- pedding
        7847 => x"00000016", -- pedding
        7848 => x"00000016", -- pedding
        7849 => x"00000016", -- pedding
        7850 => x"00000016", -- pedding
        7851 => x"00000016", -- pedding
        7852 => x"00000016", -- pedding
        7853 => x"00000016", -- pedding
        7854 => x"00000016", -- pedding
        7855 => x"00000016", -- pedding
        7856 => x"00000016", -- pedding
        7857 => x"00000016", -- pedding
        7858 => x"00000016", -- pedding
        7859 => x"00000016", -- pedding
        7860 => x"00000016", -- pedding
        7861 => x"00000016", -- pedding
        7862 => x"00000016", -- pedding
        7863 => x"00000016", -- pedding
        7864 => x"00000016", -- pedding
        7865 => x"00000016", -- pedding
        7866 => x"00000016", -- pedding
        7867 => x"00000016", -- pedding
        7868 => x"00000016", -- pedding
        7869 => x"00000016", -- pedding
        7870 => x"00000016", -- pedding
        7871 => x"00000016", -- pedding
        7872 => x"00000016", -- pedding
        7873 => x"00000016", -- pedding
        7874 => x"00000016", -- pedding
        7875 => x"00000016", -- pedding
        7876 => x"00000016", -- pedding
        7877 => x"00000016", -- pedding
        7878 => x"00000016", -- pedding
        7879 => x"00000016", -- pedding
        7880 => x"00000016", -- pedding
        7881 => x"00000016", -- pedding
        7882 => x"00000016", -- pedding
        7883 => x"00000016", -- pedding
        7884 => x"00000016", -- pedding
        7885 => x"00000016", -- pedding
        7886 => x"00000016", -- pedding
        7887 => x"00000016", -- pedding
        7888 => x"00000016", -- pedding
        7889 => x"00000016", -- pedding
        7890 => x"00000016", -- pedding
        7891 => x"00000016", -- pedding
        7892 => x"00000016", -- pedding
        7893 => x"00000016", -- pedding
        7894 => x"00000016", -- pedding
        7895 => x"00000016", -- pedding
        7896 => x"00000016", -- pedding
        7897 => x"00000016", -- pedding
        7898 => x"00000016", -- pedding
        7899 => x"00000016", -- pedding
        7900 => x"00000016", -- pedding
        7901 => x"00000016", -- pedding
        7902 => x"00000016", -- pedding
        7903 => x"00000016", -- pedding
        7904 => x"00000016", -- pedding
        7905 => x"00000016", -- pedding
        7906 => x"00000016", -- pedding
        7907 => x"00000016", -- pedding
        7908 => x"00000016", -- pedding
        7909 => x"00000016", -- pedding
        7910 => x"00000016", -- pedding
        7911 => x"00000016", -- pedding
        7912 => x"00000016", -- pedding
        7913 => x"00000016", -- pedding
        7914 => x"00000016", -- pedding
        7915 => x"00000016", -- pedding
        7916 => x"00000016", -- pedding
        7917 => x"00000016", -- pedding
        7918 => x"00000016", -- pedding
        7919 => x"00000016", -- pedding
        7920 => x"00000016", -- pedding
        7921 => x"00000016", -- pedding
        7922 => x"00000016", -- pedding
        7923 => x"00000016", -- pedding
        7924 => x"00000016", -- pedding
        7925 => x"00000016", -- pedding
        7926 => x"00000016", -- pedding
        7927 => x"00000016", -- pedding
        7928 => x"00000016", -- pedding
        7929 => x"00000016", -- pedding
        7930 => x"00000016", -- pedding
        7931 => x"00000016", -- pedding
        7932 => x"00000016", -- pedding
        7933 => x"00000016", -- pedding
        7934 => x"00000016", -- pedding
        7935 => x"00000016", -- pedding
        7936 => x"00000016", -- pedding
        7937 => x"00000016", -- pedding
        7938 => x"00000016", -- pedding
        7939 => x"00000016", -- pedding
        7940 => x"00000016", -- pedding
        7941 => x"00000016", -- pedding
        7942 => x"00000016", -- pedding
        7943 => x"00000016", -- pedding
        7944 => x"00000016", -- pedding
        7945 => x"00000016", -- pedding
        7946 => x"00000016", -- pedding
        7947 => x"00000016", -- pedding
        7948 => x"00000016", -- pedding
        7949 => x"00000016", -- pedding
        7950 => x"00000016", -- pedding
        7951 => x"00000016", -- pedding
        7952 => x"00000016", -- pedding
        7953 => x"00000016", -- pedding
        7954 => x"00000016", -- pedding
        7955 => x"00000016", -- pedding
        7956 => x"00000016", -- pedding
        7957 => x"00000016", -- pedding
        7958 => x"00000016", -- pedding
        7959 => x"00000016", -- pedding
        7960 => x"00000016", -- pedding
        7961 => x"00000016", -- pedding
        7962 => x"00000016", -- pedding
        7963 => x"00000016", -- pedding
        7964 => x"00000016", -- pedding
        7965 => x"00000016", -- pedding
        7966 => x"00000016", -- pedding
        7967 => x"00000016", -- pedding
        7968 => x"00000016", -- pedding
        7969 => x"00000016", -- pedding
        7970 => x"00000016", -- pedding
        7971 => x"00000016", -- pedding
        7972 => x"00000016", -- pedding
        7973 => x"00000016", -- pedding
        7974 => x"00000016", -- pedding
        7975 => x"00000016", -- pedding
        7976 => x"00000016", -- pedding
        7977 => x"00000016", -- pedding
        7978 => x"00000016", -- pedding
        7979 => x"00000016", -- pedding
        7980 => x"00000016", -- pedding
        7981 => x"00000016", -- pedding
        7982 => x"00000016", -- pedding
        7983 => x"00000016", -- pedding
        7984 => x"00000016", -- pedding
        7985 => x"00000016", -- pedding
        7986 => x"00000016", -- pedding
        7987 => x"00000016", -- pedding
        7988 => x"00000016", -- pedding
        7989 => x"00000016", -- pedding
        7990 => x"00000016", -- pedding
        7991 => x"00000016", -- pedding
        7992 => x"00000016", -- pedding
        7993 => x"00000016", -- pedding
        7994 => x"00000016", -- pedding
        7995 => x"00000016", -- pedding
        7996 => x"00000016", -- pedding
        7997 => x"00000016", -- pedding
        7998 => x"00000016", -- pedding
        7999 => x"00000016", -- pedding
        8000 => x"00000016", -- pedding
        8001 => x"00000016", -- pedding
        8002 => x"00000016", -- pedding
        8003 => x"00000016", -- pedding
        8004 => x"00000016", -- pedding
        8005 => x"00000016", -- pedding
        8006 => x"00000016", -- pedding
        8007 => x"00000016", -- pedding
        8008 => x"00000016", -- pedding
        8009 => x"00000016", -- pedding
        8010 => x"00000016", -- pedding
        8011 => x"00000016", -- pedding
        8012 => x"00000016", -- pedding
        8013 => x"00000016", -- pedding
        8014 => x"00000016", -- pedding
        8015 => x"00000016", -- pedding
        8016 => x"00000016", -- pedding
        8017 => x"00000016", -- pedding
        8018 => x"00000016", -- pedding
        8019 => x"00000016", -- pedding
        8020 => x"00000016", -- pedding
        8021 => x"00000016", -- pedding
        8022 => x"00000016", -- pedding
        8023 => x"00000016", -- pedding
        8024 => x"00000016", -- pedding
        8025 => x"00000016", -- pedding
        8026 => x"00000016", -- pedding
        8027 => x"00000016", -- pedding
        8028 => x"00000016", -- pedding
        8029 => x"00000016", -- pedding
        8030 => x"00000016", -- pedding
        8031 => x"00000016", -- pedding
        8032 => x"00000016", -- pedding
        8033 => x"00000016", -- pedding
        8034 => x"00000016", -- pedding
        8035 => x"00000016", -- pedding
        8036 => x"00000016", -- pedding
        8037 => x"00000016", -- pedding
        8038 => x"00000016", -- pedding
        8039 => x"00000016", -- pedding
        8040 => x"00000016", -- pedding
        8041 => x"00000016", -- pedding
        8042 => x"00000016", -- pedding
        8043 => x"00000016", -- pedding
        8044 => x"00000016", -- pedding
        8045 => x"00000016", -- pedding
        8046 => x"00000016", -- pedding
        8047 => x"00000016", -- pedding
        8048 => x"00000016", -- pedding
        8049 => x"00000016", -- pedding
        8050 => x"00000016", -- pedding
        8051 => x"00000016", -- pedding
        8052 => x"00000016", -- pedding
        8053 => x"00000016", -- pedding
        8054 => x"00000016", -- pedding
        8055 => x"00000016", -- pedding
        8056 => x"00000016", -- pedding
        8057 => x"00000016", -- pedding
        8058 => x"00000016", -- pedding
        8059 => x"00000016", -- pedding
        8060 => x"00000016", -- pedding
        8061 => x"00000016", -- pedding
        8062 => x"00000016", -- pedding
        8063 => x"00000016", -- pedding
        8064 => x"00000016", -- pedding
        8065 => x"00000016", -- pedding
        8066 => x"00000016", -- pedding
        8067 => x"00000016", -- pedding
        8068 => x"00000016", -- pedding
        8069 => x"00000016", -- pedding
        8070 => x"00000016", -- pedding
        8071 => x"00000016", -- pedding
        8072 => x"00000016", -- pedding
        8073 => x"00000016", -- pedding
        8074 => x"00000016", -- pedding
        8075 => x"00000016", -- pedding
        8076 => x"00000016", -- pedding
        8077 => x"00000016", -- pedding
        8078 => x"00000016", -- pedding
        8079 => x"00000016", -- pedding
        8080 => x"00000016", -- pedding
        8081 => x"00000016", -- pedding
        8082 => x"00000016", -- pedding
        8083 => x"00000016", -- pedding
        8084 => x"00000016", -- pedding
        8085 => x"00000016", -- pedding
        8086 => x"00000016", -- pedding
        8087 => x"00000016", -- pedding
        8088 => x"00000016", -- pedding
        8089 => x"00000016", -- pedding
        8090 => x"00000016", -- pedding
        8091 => x"00000016", -- pedding
        8092 => x"00000016", -- pedding
        8093 => x"00000016", -- pedding
        8094 => x"00000016", -- pedding
        8095 => x"00000016", -- pedding
        8096 => x"00000016", -- pedding
        8097 => x"00000016", -- pedding
        8098 => x"00000016", -- pedding
        8099 => x"00000016", -- pedding
        8100 => x"00000016", -- pedding
        8101 => x"00000016", -- pedding
        8102 => x"00000016", -- pedding
        8103 => x"00000016", -- pedding
        8104 => x"00000016", -- pedding
        8105 => x"00000016", -- pedding
        8106 => x"00000016", -- pedding
        8107 => x"00000016", -- pedding
        8108 => x"00000016", -- pedding
        8109 => x"00000016", -- pedding
        8110 => x"00000016", -- pedding
        8111 => x"00000016", -- pedding
        8112 => x"00000016", -- pedding
        8113 => x"00000016", -- pedding
        8114 => x"00000016", -- pedding
        8115 => x"00000016", -- pedding
        8116 => x"00000016", -- pedding
        8117 => x"00000016", -- pedding
        8118 => x"00000016", -- pedding
        8119 => x"00000016", -- pedding
        8120 => x"00000016", -- pedding
        8121 => x"00000016", -- pedding
        8122 => x"00000016", -- pedding
        8123 => x"00000016", -- pedding
        8124 => x"00000016", -- pedding
        8125 => x"00000016", -- pedding
        8126 => x"00000016", -- pedding
        8127 => x"00000016", -- pedding
        8128 => x"00000016", -- pedding
        8129 => x"00000016", -- pedding
        8130 => x"00000016", -- pedding
        8131 => x"00000016", -- pedding
        8132 => x"00000016", -- pedding
        8133 => x"00000016", -- pedding
        8134 => x"00000016", -- pedding
        8135 => x"00000016", -- pedding
        8136 => x"00000016", -- pedding
        8137 => x"00000016", -- pedding
        8138 => x"00000016", -- pedding
        8139 => x"00000016", -- pedding
        8140 => x"00000016", -- pedding
        8141 => x"00000016", -- pedding
        8142 => x"00000016", -- pedding
        8143 => x"00000016", -- pedding
        8144 => x"00000016", -- pedding
        8145 => x"00000016", -- pedding
        8146 => x"00000016", -- pedding
        8147 => x"00000016", -- pedding
        8148 => x"00000016", -- pedding
        8149 => x"00000016", -- pedding
        8150 => x"00000016", -- pedding
        8151 => x"00000016", -- pedding
        8152 => x"00000016", -- pedding
        8153 => x"00000016", -- pedding
        8154 => x"00000016", -- pedding
        8155 => x"00000016", -- pedding
        8156 => x"00000016", -- pedding
        8157 => x"00000016", -- pedding
        8158 => x"00000016", -- pedding
        8159 => x"00000016", -- pedding
        8160 => x"00000016", -- pedding
        8161 => x"00000016", -- pedding
        8162 => x"00000016", -- pedding
        8163 => x"00000016", -- pedding
        8164 => x"00000016", -- pedding
        8165 => x"00000016", -- pedding
        8166 => x"00000016", -- pedding
        8167 => x"00000016", -- pedding
        8168 => x"00000016", -- pedding
        8169 => x"00000016", -- pedding
        8170 => x"00000016", -- pedding
        8171 => x"00000016", -- pedding
        8172 => x"00000016", -- pedding
        8173 => x"00000016", -- pedding
        8174 => x"00000016", -- pedding
        8175 => x"00000016", -- pedding
        8176 => x"00000016", -- pedding
        8177 => x"00000016", -- pedding
        8178 => x"00000016", -- pedding
        8179 => x"00000016", -- pedding
        8180 => x"00000016", -- pedding
        8181 => x"00000016", -- pedding
        8182 => x"00000016", -- pedding
        8183 => x"00000016", -- pedding
        8184 => x"00000016", -- pedding
        8185 => x"00000016", -- pedding
        8186 => x"00000016", -- pedding
        8187 => x"00000016", -- pedding
        8188 => x"00000016", -- pedding
        8189 => x"00000016", -- pedding
        8190 => x"00000016", -- pedding
        8191 => x"00000016", -- pedding


others => x"00000000"
	);


begin

	process(i_clk)
	begin
		if rising_edge(i_clk) then
			-- memory write --
			if i_we = '1' then
				mem(to_integer(unsigned(i_w_addr))) <= i_data;
			end if;
			-- memory read --
			o_data <= mem(to_integer(unsigned(i_r_addr)));

		end if;
	end process;

end architecture arch;