
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity ram is
	generic
	(
		DATA_WIDTH : natural := 32;		    -- 4 byte one line of memory
		ADDR_WIDTH : natural := 13			    -- 24576 bytes size of memory
	);

	port(
		i_clk    : in  std_logic;
		i_r_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		i_data   : in  std_logic_vector(DATA_WIDTH-1 downto 0);
		i_we     : in  std_logic;
		i_w_addr : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
		o_data   : out std_logic_vector(DATA_WIDTH-1 downto 0)
	);
end entity ram;

architecture arch of ram is

	type ram_t is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(DATA_WIDTH-1 downto 0);


-- GENERATED BY BC_MEM_PACKER

-- DATE: Thu May 18 16:01:02 2017

	signal mem : ram_t := (

--			***** COLOR PALLETE *****

		-- fellas
		0 =>	x"000C4CC8",
		1 =>	x"00A8D8FC",
		2 =>	x"00000000",
		3 =>	x"00EC3820",
		4 =>	x"0000A800",
		5 =>	x"00FCFCFC",
		6 =>	x"00747474",
		7 =>	x"00C0C0C0",
--      Link colors
        8 =>    x"00303030",
        9 =>    x"000CCB83",
        10 =>   x"002C98D8",
        11 =>   x"00004B7B",
        12 =>   x"00FFD9D9",
        13 =>   x"00003299",
        14 =>   x"00B1DFF8",
        15 =>   x"00FFFFFF",
        16 =>   x"008E0018",
        17 =>   x"00FF898E",
        18 =>   x"00000000",
        19 =>   x"00006E8A",
        20 =>   x"00002E55",
        21 =>   x"00CBC74D",
        22 =>   x"00E32F47",
        23 =>   x"00173B00",
        24 =>   x"00007A3E",
        25 =>   x"007ED14A",
        26 =>   x"0000311D",
        27 =>   x"0000675B",
        28 =>   x"000AB4B9",
        29 =>   x"00003D00",
        30 =>   x"00008200",
        31 =>   x"003FD65B",
        32 =>   x"00656565",
        33 =>   x"00B9B9B9",
        34 =>   x"00AFAFAF",
-- 		enemie colors
		35 =>	x"00c0c0c0",
		36 => 	x"000038f8",
		37 => 	x"00bc0000",
		38 =>	x"00ff8868",
		39 => 	x"00ffffff",
																															-- map colors
																															40 => x"00000000",
																															41 => x"00120a00",
																															42 => x"00513800",
																															43 => x"00735200",
																															44 => x"007f5b00",
																															45 => x"007e5a00",
																															46 => x"00523900",
																															47 => x"00271900",
																															48 => x"00080400",
																															49 => x"00010000",
																															50 => x"00d8e800",
																															51 => x"00000a00",
																															52 => x"0000d600",
																															53 => x"00020202",
																															54 => x"00010101",
																															55 => x"00010100",
																															56 => x"00030600",
																															57 => x"00105ce4",
																															58 => x"0044a0fc",
																															59 => x"00bc0000",
																															60 => x"005800e4",
																															61 => x"00020100",
																															62 => x"00f85800",
		63 =>	x"003199FF", -- Unused

            --  ADDED SPRITES HERE
          -- RUPEE SPRITE
		64 => x"0202020F",
		65 => x"3C020202",
		66 => x"02020202",
		67 => x"02020202",
		68 => x"02020F0F",
		69 => x"3C3C0202",
		70 => x"02020202",
		71 => x"02020202",
		72 => x"020F0F0F",
		73 => x"3C3C3C02",
		74 => x"02020202",
		75 => x"02020202",
		76 => x"0F3C0F3C",
		77 => x"023C023C",
		78 => x"02020202",
		79 => x"02020202",
		80 => x"0F0F3C3C",
		81 => x"3C023C3C",
		82 => x"02020202",
		83 => x"02020202",
		84 => x"0F0F3C3C",
		85 => x"3C023C3C",
		86 => x"02020202",
		87 => x"02020202",
		88 => x"0F0F3C3C",
		89 => x"3C023C3C",
		90 => x"02020202",
		91 => x"02020202",
		92 => x"0F0F3C3C",
		93 => x"3C023C3C",
		94 => x"02020202",
		95 => x"02020202",
		96 => x"0F0F3C3C",
		97 => x"3C023C3C",
		98 => x"02020202",
		99 => x"02020202",
		100 => x"0F0F3C3C",
		101 => x"3C023C3C",
		102 => x"02020202",
		103 => x"02020202",
		104 => x"0F0F3C3C",
		105 => x"3C023C3C",
		106 => x"02020202",
		107 => x"02020202",
		108 => x"0F3C0F3C",
		109 => x"3C023C3C",
		110 => x"02020202",
		111 => x"02020202",
		112 => x"3C3C3C0F",
		113 => x"023C023C",
		114 => x"02020202",
		115 => x"02020202",
		116 => x"023C3C3C",
		117 => x"3C3C3C02",
		118 => x"02020202",
		119 => x"02020202",
		120 => x"02023C3C",
		121 => x"3C3C0202",
		122 => x"02020202",
		123 => x"02020202",
		124 => x"0202023C",
		125 => x"3C020202",
		126 => x"02020202",
		127 => x"02020202",

          -- BOMB SPRITE
		128 => x"02020202",
		129 => x"020F0202",
		130 => x"02020202",
		131 => x"02020202",
		132 => x"02020202",
		133 => x"020F0202",
		134 => x"02020202",
		135 => x"02020202",
		136 => x"02020202",
		137 => x"02020F02",
		138 => x"02020202",
		139 => x"02020202",
		140 => x"02020202",
		141 => x"0202020F",
		142 => x"02020202",
		143 => x"02020202",
		144 => x"02020202",
		145 => x"0202020F",
		146 => x"02020202",
		147 => x"02020202",
		148 => x"02020202",
		149 => x"02020F02",
		150 => x"02020202",
		151 => x"02020202",
		152 => x"02020D0D",
		153 => x"0D0D0202",
		154 => x"02020202",
		155 => x"02020202",
		156 => x"020D2E2E",
		157 => x"0D0D0D02",
		158 => x"02020202",
		159 => x"02020202",
		160 => x"0D2E0F2E",
		161 => x"0D0D0D0D",
		162 => x"02020202",
		163 => x"02020202",
		164 => x"0D2E2E0D",
		165 => x"0D0D0D0D",
		166 => x"02020202",
		167 => x"02020202",
		168 => x"0D0D0D0D",
		169 => x"0D0D0D0D",
		170 => x"02020202",
		171 => x"02020202",
		172 => x"0D0D0D0D",
		173 => x"0D0D0D0D",
		174 => x"02020202",
		175 => x"02020202",
		176 => x"020D0D0D",
		177 => x"0D0D0D02",
		178 => x"02020202",
		179 => x"02020202",
		180 => x"02020D0D",
		181 => x"0D0D0202",
		182 => x"02020202",
		183 => x"02020202",
		184 => x"02020202",
		185 => x"02020202",
		186 => x"02020202",
		187 => x"02020202",
		188 => x"02020202",
		189 => x"02020202",
		190 => x"02020202",
		191 => x"02020202",

--			***** 16x16 IMAGES *****
--			OVERWORLD SPRITES

      --  sprite 0

			                --  sprite 0
			        255 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        256 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        257 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        258 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        259 => x"00000000",		-- colors: 40, 40, 40, 40
			        260 => x"00000000",		-- colors: 40, 40, 40, 40
			        261 => x"00000000",		-- colors: 40, 40, 40, 40
			        262 => x"00000000",		-- colors: 40, 40, 40, 40
			        263 => x"00000000",		-- colors: 40, 40, 40, 40
			        264 => x"00000000",		-- colors: 40, 40, 40, 40
			        265 => x"00000000",		-- colors: 40, 40, 40, 40
			        266 => x"00000000",		-- colors: 40, 40, 40, 40
			        267 => x"00000000",		-- colors: 40, 40, 40, 40
			        268 => x"00000000",		-- colors: 40, 40, 40, 40
			        269 => x"00000000",		-- colors: 40, 40, 40, 40
			        270 => x"00000000",		-- colors: 40, 40, 40, 40
			        271 => x"00000000",		-- colors: 40, 40, 40, 40
			        272 => x"00000000",		-- colors: 40, 40, 40, 40
			        273 => x"00000000",		-- colors: 40, 40, 40, 40
			        274 => x"00000000",		-- colors: 40, 40, 40, 40
			        275 => x"00000000",		-- colors: 40, 40, 40, 40
			        276 => x"00000000",		-- colors: 40, 40, 40, 40
			        277 => x"00000000",		-- colors: 40, 40, 40, 40
			        278 => x"00000000",		-- colors: 40, 40, 40, 40
			        279 => x"00000000",		-- colors: 40, 40, 40, 40
			        280 => x"00000000",		-- colors: 40, 40, 40, 40
			        281 => x"00000000",		-- colors: 40, 40, 40, 40
			        282 => x"00000000",		-- colors: 40, 40, 40, 40
			        283 => x"00000000",		-- colors: 40, 40, 40, 40
			        284 => x"00000000",		-- colors: 40, 40, 40, 40
			        285 => x"00000000",		-- colors: 40, 40, 40, 40
			        286 => x"00000000",		-- colors: 40, 40, 40, 40
			        287 => x"00000000",		-- colors: 40, 40, 40, 40
			        288 => x"00000000",		-- colors: 40, 40, 40, 40
			        289 => x"00000000",		-- colors: 40, 40, 40, 40
			        290 => x"00000000",		-- colors: 40, 40, 40, 40
			        291 => x"00000000",		-- colors: 40, 40, 40, 40
			        292 => x"00000000",		-- colors: 40, 40, 40, 40
			        293 => x"00000000",		-- colors: 40, 40, 40, 40
			        294 => x"00000000",		-- colors: 40, 40, 40, 40
			        295 => x"00000000",		-- colors: 40, 40, 40, 40
			        296 => x"00000000",		-- colors: 40, 40, 40, 40
			        297 => x"00000000",		-- colors: 40, 40, 40, 40
			        298 => x"00000000",		-- colors: 40, 40, 40, 40
			        299 => x"00000000",		-- colors: 40, 40, 40, 40
			        300 => x"00000000",		-- colors: 40, 40, 40, 40
			        301 => x"00000000",		-- colors: 40, 40, 40, 40
			        302 => x"00000000",		-- colors: 40, 40, 40, 40
			        303 => x"00000000",		-- colors: 40, 40, 40, 40
			        304 => x"00000000",		-- colors: 40, 40, 40, 40
			        305 => x"00000000",		-- colors: 40, 40, 40, 40
			        306 => x"00000000",		-- colors: 40, 40, 40, 40
			        307 => x"00000000",		-- colors: 40, 40, 40, 40
			        308 => x"00000000",		-- colors: 40, 40, 40, 40
			        309 => x"00000000",		-- colors: 40, 40, 40, 40
			        310 => x"00000000",		-- colors: 40, 40, 40, 40
			        311 => x"00000000",		-- colors: 40, 40, 40, 40
			        312 => x"00000000",		-- colors: 40, 40, 40, 40
			        313 => x"00000000",		-- colors: 40, 40, 40, 40
			        314 => x"00000000",		-- colors: 40, 40, 40, 40
			        315 => x"00000000",		-- colors: 40, 40, 40, 40
			        316 => x"00000000",		-- colors: 40, 40, 40, 40
			        317 => x"00000000",		-- colors: 40, 40, 40, 40
			        318 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 1
			        319 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        320 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        321 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        322 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        323 => x"00000000",		-- colors: 40, 40, 40, 40
			        324 => x"00000000",		-- colors: 40, 40, 40, 40
			        325 => x"00000000",		-- colors: 40, 40, 40, 40
			        326 => x"00000000",		-- colors: 40, 40, 40, 40
			        327 => x"00000000",		-- colors: 40, 40, 40, 40
			        328 => x"00000000",		-- colors: 40, 40, 40, 40
			        329 => x"00000000",		-- colors: 40, 40, 40, 40
			        330 => x"00000000",		-- colors: 40, 40, 40, 40
			        331 => x"00000000",		-- colors: 40, 40, 40, 40
			        332 => x"00000000",		-- colors: 40, 40, 40, 40
			        333 => x"00000000",		-- colors: 40, 40, 40, 40
			        334 => x"00000000",		-- colors: 40, 40, 40, 40
			        335 => x"00000000",		-- colors: 40, 40, 40, 40
			        336 => x"00000000",		-- colors: 40, 40, 40, 40
			        337 => x"00000000",		-- colors: 40, 40, 40, 40
			        338 => x"00000000",		-- colors: 40, 40, 40, 40
			        339 => x"00000000",		-- colors: 40, 40, 40, 40
			        340 => x"00000000",		-- colors: 40, 40, 40, 40
			        341 => x"00000000",		-- colors: 40, 40, 40, 40
			        342 => x"00000000",		-- colors: 40, 40, 40, 40
			        343 => x"00000000",		-- colors: 40, 40, 40, 40
			        344 => x"00000000",		-- colors: 40, 40, 40, 40
			        345 => x"00000000",		-- colors: 40, 40, 40, 40
			        346 => x"00000000",		-- colors: 40, 40, 40, 40
			        347 => x"00000000",		-- colors: 40, 40, 40, 40
			        348 => x"00000000",		-- colors: 40, 40, 40, 40
			        349 => x"00000000",		-- colors: 40, 40, 40, 40
			        350 => x"00000000",		-- colors: 40, 40, 40, 40
			        351 => x"00000000",		-- colors: 40, 40, 40, 40
			        352 => x"00000000",		-- colors: 40, 40, 40, 40
			        353 => x"00000000",		-- colors: 40, 40, 40, 40
			        354 => x"00000000",		-- colors: 40, 40, 40, 40
			        355 => x"00000000",		-- colors: 40, 40, 40, 40
			        356 => x"00000000",		-- colors: 40, 40, 40, 40
			        357 => x"00000000",		-- colors: 40, 40, 40, 40
			        358 => x"00000000",		-- colors: 40, 40, 40, 40
			        359 => x"00000000",		-- colors: 40, 40, 40, 40
			        360 => x"00000000",		-- colors: 40, 40, 40, 40
			        361 => x"00000000",		-- colors: 40, 40, 40, 40
			        362 => x"00000000",		-- colors: 40, 40, 40, 40
			        363 => x"00000000",		-- colors: 40, 40, 40, 40
			        364 => x"00000000",		-- colors: 40, 40, 40, 40
			        365 => x"00000000",		-- colors: 40, 40, 40, 40
			        366 => x"00000000",		-- colors: 40, 40, 40, 40
			        367 => x"00000000",		-- colors: 40, 40, 40, 40
			        368 => x"00000000",		-- colors: 40, 40, 40, 40
			        369 => x"00000000",		-- colors: 40, 40, 40, 40
			        370 => x"00000000",		-- colors: 40, 40, 40, 40
			        371 => x"00000000",		-- colors: 40, 40, 40, 40
			        372 => x"00000000",		-- colors: 40, 40, 40, 40
			        373 => x"00000000",		-- colors: 40, 40, 40, 40
			        374 => x"00000000",		-- colors: 40, 40, 40, 40
			        375 => x"00000000",		-- colors: 40, 40, 40, 40
			        376 => x"00000000",		-- colors: 40, 40, 40, 40
			        377 => x"00000000",		-- colors: 40, 40, 40, 40
			        378 => x"00000000",		-- colors: 40, 40, 40, 40
			        379 => x"00000000",		-- colors: 40, 40, 40, 40
			        380 => x"00000000",		-- colors: 40, 40, 40, 40
			        381 => x"00000000",		-- colors: 40, 40, 40, 40
			        382 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 2
			        383 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        384 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        385 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        386 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        387 => x"00000000",		-- colors: 40, 40, 40, 40
			        388 => x"00000000",		-- colors: 40, 40, 40, 40
			        389 => x"00000000",		-- colors: 40, 40, 40, 40
			        390 => x"00000000",		-- colors: 40, 40, 40, 40
			        391 => x"00000000",		-- colors: 40, 40, 40, 40
			        392 => x"00000000",		-- colors: 40, 40, 40, 40
			        393 => x"00000000",		-- colors: 40, 40, 40, 40
			        394 => x"00000000",		-- colors: 40, 40, 40, 40
			        395 => x"00000000",		-- colors: 40, 40, 40, 40
			        396 => x"00000000",		-- colors: 40, 40, 40, 40
			        397 => x"00000000",		-- colors: 40, 40, 40, 40
			        398 => x"00000000",		-- colors: 40, 40, 40, 40
			        399 => x"00000000",		-- colors: 40, 40, 40, 40
			        400 => x"00000000",		-- colors: 40, 40, 40, 40
			        401 => x"00000000",		-- colors: 40, 40, 40, 40
			        402 => x"00000000",		-- colors: 40, 40, 40, 40
			        403 => x"00000000",		-- colors: 40, 40, 40, 40
			        404 => x"00000000",		-- colors: 40, 40, 40, 40
			        405 => x"00000000",		-- colors: 40, 40, 40, 40
			        406 => x"00000000",		-- colors: 40, 40, 40, 40
			        407 => x"00000000",		-- colors: 40, 40, 40, 40
			        408 => x"00000000",		-- colors: 40, 40, 40, 40
			        409 => x"00000000",		-- colors: 40, 40, 40, 40
			        410 => x"00000000",		-- colors: 40, 40, 40, 40
			        411 => x"00000000",		-- colors: 40, 40, 40, 40
			        412 => x"00000000",		-- colors: 40, 40, 40, 40
			        413 => x"00000000",		-- colors: 40, 40, 40, 40
			        414 => x"00000000",		-- colors: 40, 40, 40, 40
			        415 => x"00000000",		-- colors: 40, 40, 40, 40
			        416 => x"00000000",		-- colors: 40, 40, 40, 40
			        417 => x"00000000",		-- colors: 40, 40, 40, 40
			        418 => x"00000000",		-- colors: 40, 40, 40, 40
			        419 => x"00000000",		-- colors: 40, 40, 40, 40
			        420 => x"00000000",		-- colors: 40, 40, 40, 40
			        421 => x"00000000",		-- colors: 40, 40, 40, 40
			        422 => x"00000000",		-- colors: 40, 40, 40, 40
			        423 => x"00000000",		-- colors: 40, 40, 40, 40
			        424 => x"00000000",		-- colors: 40, 40, 40, 40
			        425 => x"00000000",		-- colors: 40, 40, 40, 40
			        426 => x"00000000",		-- colors: 40, 40, 40, 40
			        427 => x"00000000",		-- colors: 40, 40, 40, 40
			        428 => x"00000000",		-- colors: 40, 40, 40, 40
			        429 => x"00000000",		-- colors: 40, 40, 40, 40
			        430 => x"00000000",		-- colors: 40, 40, 40, 40
			        431 => x"00000000",		-- colors: 40, 40, 40, 40
			        432 => x"00000000",		-- colors: 40, 40, 40, 40
			        433 => x"00000000",		-- colors: 40, 40, 40, 40
			        434 => x"00000000",		-- colors: 40, 40, 40, 40
			        435 => x"00000000",		-- colors: 40, 40, 40, 40
			        436 => x"00000000",		-- colors: 40, 40, 40, 40
			        437 => x"00000000",		-- colors: 40, 40, 40, 40
			        438 => x"00000000",		-- colors: 40, 40, 40, 40
			        439 => x"00000000",		-- colors: 40, 40, 40, 40
			        440 => x"00000000",		-- colors: 40, 40, 40, 40
			        441 => x"00000000",		-- colors: 40, 40, 40, 40
			        442 => x"00000000",		-- colors: 40, 40, 40, 40
			        443 => x"00000000",		-- colors: 40, 40, 40, 40
			        444 => x"00000000",		-- colors: 40, 40, 40, 40
			        445 => x"00000000",		-- colors: 40, 40, 40, 40
			        446 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 3
			        447 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        448 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        449 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        450 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        451 => x"00000000",		-- colors: 40, 40, 40, 40
			        452 => x"00000000",		-- colors: 40, 40, 40, 40
			        453 => x"00000000",		-- colors: 40, 40, 40, 40
			        454 => x"00000000",		-- colors: 40, 40, 40, 40
			        455 => x"00000000",		-- colors: 40, 40, 40, 40
			        456 => x"00000000",		-- colors: 40, 40, 40, 40
			        457 => x"00000000",		-- colors: 40, 40, 40, 40
			        458 => x"00000000",		-- colors: 40, 40, 40, 40
			        459 => x"00000000",		-- colors: 40, 40, 40, 40
			        460 => x"00000000",		-- colors: 40, 40, 40, 40
			        461 => x"00000000",		-- colors: 40, 40, 40, 40
			        462 => x"00000000",		-- colors: 40, 40, 40, 40
			        463 => x"00000000",		-- colors: 40, 40, 40, 40
			        464 => x"00000000",		-- colors: 40, 40, 40, 40
			        465 => x"00000000",		-- colors: 40, 40, 40, 40
			        466 => x"00000000",		-- colors: 40, 40, 40, 40
			        467 => x"00000000",		-- colors: 40, 40, 40, 40
			        468 => x"00000000",		-- colors: 40, 40, 40, 40
			        469 => x"00000000",		-- colors: 40, 40, 40, 40
			        470 => x"00000000",		-- colors: 40, 40, 40, 40
			        471 => x"00000000",		-- colors: 40, 40, 40, 40
			        472 => x"00000000",		-- colors: 40, 40, 40, 40
			        473 => x"00000000",		-- colors: 40, 40, 40, 40
			        474 => x"00000000",		-- colors: 40, 40, 40, 40
			        475 => x"00000000",		-- colors: 40, 40, 40, 40
			        476 => x"00000000",		-- colors: 40, 40, 40, 40
			        477 => x"00000000",		-- colors: 40, 40, 40, 40
			        478 => x"00000000",		-- colors: 40, 40, 40, 40
			        479 => x"00000000",		-- colors: 40, 40, 40, 40
			        480 => x"00000000",		-- colors: 40, 40, 40, 40
			        481 => x"00000000",		-- colors: 40, 40, 40, 40
			        482 => x"00000000",		-- colors: 40, 40, 40, 40
			        483 => x"00000000",		-- colors: 40, 40, 40, 40
			        484 => x"00000000",		-- colors: 40, 40, 40, 40
			        485 => x"00000000",		-- colors: 40, 40, 40, 40
			        486 => x"00000000",		-- colors: 40, 40, 40, 40
			        487 => x"00000000",		-- colors: 40, 40, 40, 40
			        488 => x"00000000",		-- colors: 40, 40, 40, 40
			        489 => x"00000000",		-- colors: 40, 40, 40, 40
			        490 => x"00000000",		-- colors: 40, 40, 40, 40
			        491 => x"00000000",		-- colors: 40, 40, 40, 40
			        492 => x"00000000",		-- colors: 40, 40, 40, 40
			        493 => x"00000000",		-- colors: 40, 40, 40, 40
			        494 => x"00000000",		-- colors: 40, 40, 40, 40
			        495 => x"00000000",		-- colors: 40, 40, 40, 40
			        496 => x"00000000",		-- colors: 40, 40, 40, 40
			        497 => x"00000000",		-- colors: 40, 40, 40, 40
			        498 => x"00000000",		-- colors: 40, 40, 40, 40
			        499 => x"00000000",		-- colors: 40, 40, 40, 40
			        500 => x"00000000",		-- colors: 40, 40, 40, 40
			        501 => x"00000000",		-- colors: 40, 40, 40, 40
			        502 => x"00000000",		-- colors: 40, 40, 40, 40
			        503 => x"00000000",		-- colors: 40, 40, 40, 40
			        504 => x"00000000",		-- colors: 40, 40, 40, 40
			        505 => x"00000000",		-- colors: 40, 40, 40, 40
			        506 => x"00000000",		-- colors: 40, 40, 40, 40
			        507 => x"00000000",		-- colors: 40, 40, 40, 40
			        508 => x"00000000",		-- colors: 40, 40, 40, 40
			        509 => x"00000000",		-- colors: 40, 40, 40, 40
			        510 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 4
			        511 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        512 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        513 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        514 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        515 => x"00000000",		-- colors: 40, 40, 40, 40
			        516 => x"00000000",		-- colors: 40, 40, 40, 40
			        517 => x"00000000",		-- colors: 40, 40, 40, 40
			        518 => x"00000000",		-- colors: 40, 40, 40, 40
			        519 => x"00000000",		-- colors: 40, 40, 40, 40
			        520 => x"00000000",		-- colors: 40, 40, 40, 40
			        521 => x"00000000",		-- colors: 40, 40, 40, 40
			        522 => x"00000000",		-- colors: 40, 40, 40, 40
			        523 => x"00000000",		-- colors: 40, 40, 40, 40
			        524 => x"00000000",		-- colors: 40, 40, 40, 40
			        525 => x"00000000",		-- colors: 40, 40, 40, 40
			        526 => x"00000000",		-- colors: 40, 40, 40, 40
			        527 => x"00000000",		-- colors: 40, 40, 40, 40
			        528 => x"00000000",		-- colors: 40, 40, 40, 40
			        529 => x"00000000",		-- colors: 40, 40, 40, 40
			        530 => x"00000000",		-- colors: 40, 40, 40, 40
			        531 => x"00000000",		-- colors: 40, 40, 40, 40
			        532 => x"00000000",		-- colors: 40, 40, 40, 40
			        533 => x"00000000",		-- colors: 40, 40, 40, 40
			        534 => x"00000000",		-- colors: 40, 40, 40, 40
			        535 => x"00000000",		-- colors: 40, 40, 40, 40
			        536 => x"00000000",		-- colors: 40, 40, 40, 40
			        537 => x"00000000",		-- colors: 40, 40, 40, 40
			        538 => x"00000000",		-- colors: 40, 40, 40, 40
			        539 => x"00000000",		-- colors: 40, 40, 40, 40
			        540 => x"00000000",		-- colors: 40, 40, 40, 40
			        541 => x"00000000",		-- colors: 40, 40, 40, 40
			        542 => x"00000000",		-- colors: 40, 40, 40, 40
			        543 => x"00000000",		-- colors: 40, 40, 40, 40
			        544 => x"00000000",		-- colors: 40, 40, 40, 40
			        545 => x"00000000",		-- colors: 40, 40, 40, 40
			        546 => x"00000000",		-- colors: 40, 40, 40, 40
			        547 => x"00000000",		-- colors: 40, 40, 40, 40
			        548 => x"00000000",		-- colors: 40, 40, 40, 40
			        549 => x"00000000",		-- colors: 40, 40, 40, 40
			        550 => x"00000000",		-- colors: 40, 40, 40, 40
			        551 => x"00000000",		-- colors: 40, 40, 40, 40
			        552 => x"00000000",		-- colors: 40, 40, 40, 40
			        553 => x"00000000",		-- colors: 40, 40, 40, 40
			        554 => x"00000000",		-- colors: 40, 40, 40, 40
			        555 => x"00000000",		-- colors: 40, 40, 40, 40
			        556 => x"00000000",		-- colors: 40, 40, 40, 40
			        557 => x"00000000",		-- colors: 40, 40, 40, 40
			        558 => x"00000000",		-- colors: 40, 40, 40, 40
			        559 => x"00000000",		-- colors: 40, 40, 40, 40
			        560 => x"00000000",		-- colors: 40, 40, 40, 40
			        561 => x"00000000",		-- colors: 40, 40, 40, 40
			        562 => x"00000000",		-- colors: 40, 40, 40, 40
			        563 => x"00000000",		-- colors: 40, 40, 40, 40
			        564 => x"00000000",		-- colors: 40, 40, 40, 40
			        565 => x"00000000",		-- colors: 40, 40, 40, 40
			        566 => x"00000000",		-- colors: 40, 40, 40, 40
			        567 => x"00000000",		-- colors: 40, 40, 40, 40
			        568 => x"00000000",		-- colors: 40, 40, 40, 40
			        569 => x"00000000",		-- colors: 40, 40, 40, 40
			        570 => x"00000000",		-- colors: 40, 40, 40, 40
			        571 => x"00000000",		-- colors: 40, 40, 40, 40
			        572 => x"00000000",		-- colors: 40, 40, 40, 40
			        573 => x"00000000",		-- colors: 40, 40, 40, 40
			        574 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 5
			        575 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        576 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        577 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        578 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        579 => x"00000000",		-- colors: 40, 40, 40, 40
			        580 => x"00000000",		-- colors: 40, 40, 40, 40
			        581 => x"00000000",		-- colors: 40, 40, 40, 40
			        582 => x"00000000",		-- colors: 40, 40, 40, 40
			        583 => x"00000000",		-- colors: 40, 40, 40, 40
			        584 => x"00000000",		-- colors: 40, 40, 40, 40
			        585 => x"00000000",		-- colors: 40, 40, 40, 40
			        586 => x"00000000",		-- colors: 40, 40, 40, 40
			        587 => x"00000000",		-- colors: 40, 40, 40, 40
			        588 => x"00000000",		-- colors: 40, 40, 40, 40
			        589 => x"00000000",		-- colors: 40, 40, 40, 40
			        590 => x"00000000",		-- colors: 40, 40, 40, 40
			        591 => x"00000000",		-- colors: 40, 40, 40, 40
			        592 => x"00000000",		-- colors: 40, 40, 40, 40
			        593 => x"00000000",		-- colors: 40, 40, 40, 40
			        594 => x"00000000",		-- colors: 40, 40, 40, 40
			        595 => x"00000000",		-- colors: 40, 40, 40, 40
			        596 => x"00000000",		-- colors: 40, 40, 40, 40
			        597 => x"00000000",		-- colors: 40, 40, 40, 40
			        598 => x"00000000",		-- colors: 40, 40, 40, 40
			        599 => x"00000000",		-- colors: 40, 40, 40, 40
			        600 => x"00000000",		-- colors: 40, 40, 40, 40
			        601 => x"00000000",		-- colors: 40, 40, 40, 40
			        602 => x"00000000",		-- colors: 40, 40, 40, 40
			        603 => x"00000000",		-- colors: 40, 40, 40, 40
			        604 => x"00000000",		-- colors: 40, 40, 40, 40
			        605 => x"00000000",		-- colors: 40, 40, 40, 40
			        606 => x"00000000",		-- colors: 40, 40, 40, 40
			        607 => x"00000000",		-- colors: 40, 40, 40, 40
			        608 => x"00000000",		-- colors: 40, 40, 40, 40
			        609 => x"00000000",		-- colors: 40, 40, 40, 40
			        610 => x"00000000",		-- colors: 40, 40, 40, 40
			        611 => x"00000000",		-- colors: 40, 40, 40, 40
			        612 => x"00000000",		-- colors: 40, 40, 40, 40
			        613 => x"00000000",		-- colors: 40, 40, 40, 40
			        614 => x"00000000",		-- colors: 40, 40, 40, 40
			        615 => x"00000000",		-- colors: 40, 40, 40, 40
			        616 => x"00000000",		-- colors: 40, 40, 40, 40
			        617 => x"00000000",		-- colors: 40, 40, 40, 40
			        618 => x"00000000",		-- colors: 40, 40, 40, 40
			        619 => x"00000000",		-- colors: 40, 40, 40, 40
			        620 => x"00000000",		-- colors: 40, 40, 40, 40
			        621 => x"00000000",		-- colors: 40, 40, 40, 40
			        622 => x"00000000",		-- colors: 40, 40, 40, 40
			        623 => x"00000000",		-- colors: 40, 40, 40, 40
			        624 => x"00000000",		-- colors: 40, 40, 40, 40
			        625 => x"00000000",		-- colors: 40, 40, 40, 40
			        626 => x"00000000",		-- colors: 40, 40, 40, 40
			        627 => x"00000000",		-- colors: 40, 40, 40, 40
			        628 => x"00000000",		-- colors: 40, 40, 40, 40
			        629 => x"00000000",		-- colors: 40, 40, 40, 40
			        630 => x"00000000",		-- colors: 40, 40, 40, 40
			        631 => x"00000000",		-- colors: 40, 40, 40, 40
			        632 => x"00000000",		-- colors: 40, 40, 40, 40
			        633 => x"00000000",		-- colors: 40, 40, 40, 40
			        634 => x"00000000",		-- colors: 40, 40, 40, 40
			        635 => x"00000000",		-- colors: 40, 40, 40, 40
			        636 => x"00000000",		-- colors: 40, 40, 40, 40
			        637 => x"00000000",		-- colors: 40, 40, 40, 40
			        638 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 6
			        639 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        640 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        641 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        642 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        643 => x"00000000",		-- colors: 40, 40, 40, 40
			        644 => x"00000000",		-- colors: 40, 40, 40, 40
			        645 => x"00000000",		-- colors: 40, 40, 40, 40
			        646 => x"00000000",		-- colors: 40, 40, 40, 40
			        647 => x"00000000",		-- colors: 40, 40, 40, 40
			        648 => x"00000000",		-- colors: 40, 40, 40, 40
			        649 => x"00000000",		-- colors: 40, 40, 40, 40
			        650 => x"00000000",		-- colors: 40, 40, 40, 40
			        651 => x"00000000",		-- colors: 40, 40, 40, 40
			        652 => x"00000000",		-- colors: 40, 40, 40, 40
			        653 => x"00000000",		-- colors: 40, 40, 40, 40
			        654 => x"00000000",		-- colors: 40, 40, 40, 40
			        655 => x"00000000",		-- colors: 40, 40, 40, 40
			        656 => x"00000000",		-- colors: 40, 40, 40, 40
			        657 => x"00000000",		-- colors: 40, 40, 40, 40
			        658 => x"00000000",		-- colors: 40, 40, 40, 40
			        659 => x"00000000",		-- colors: 40, 40, 40, 40
			        660 => x"00000000",		-- colors: 40, 40, 40, 40
			        661 => x"00000000",		-- colors: 40, 40, 40, 40
			        662 => x"00000000",		-- colors: 40, 40, 40, 40
			        663 => x"00000000",		-- colors: 40, 40, 40, 40
			        664 => x"00000000",		-- colors: 40, 40, 40, 40
			        665 => x"00000000",		-- colors: 40, 40, 40, 40
			        666 => x"00000000",		-- colors: 40, 40, 40, 40
			        667 => x"00000000",		-- colors: 40, 40, 40, 40
			        668 => x"00000000",		-- colors: 40, 40, 40, 40
			        669 => x"00000000",		-- colors: 40, 40, 40, 40
			        670 => x"00000000",		-- colors: 40, 40, 40, 40
			        671 => x"00000000",		-- colors: 40, 40, 40, 40
			        672 => x"00000000",		-- colors: 40, 40, 40, 40
			        673 => x"00000000",		-- colors: 40, 40, 40, 40
			        674 => x"00000000",		-- colors: 40, 40, 40, 40
			        675 => x"00000000",		-- colors: 40, 40, 40, 40
			        676 => x"00000000",		-- colors: 40, 40, 40, 40
			        677 => x"00000000",		-- colors: 40, 40, 40, 40
			        678 => x"00000000",		-- colors: 40, 40, 40, 40
			        679 => x"00000000",		-- colors: 40, 40, 40, 40
			        680 => x"00000000",		-- colors: 40, 40, 40, 40
			        681 => x"00000000",		-- colors: 40, 40, 40, 40
			        682 => x"00000000",		-- colors: 40, 40, 40, 40
			        683 => x"00000000",		-- colors: 40, 40, 40, 40
			        684 => x"00000000",		-- colors: 40, 40, 40, 40
			        685 => x"00000000",		-- colors: 40, 40, 40, 40
			        686 => x"00000000",		-- colors: 40, 40, 40, 40
			        687 => x"00000000",		-- colors: 40, 40, 40, 40
			        688 => x"00000000",		-- colors: 40, 40, 40, 40
			        689 => x"00000000",		-- colors: 40, 40, 40, 40
			        690 => x"00000000",		-- colors: 40, 40, 40, 40
			        691 => x"00000000",		-- colors: 40, 40, 40, 40
			        692 => x"00000000",		-- colors: 40, 40, 40, 40
			        693 => x"00000000",		-- colors: 40, 40, 40, 40
			        694 => x"00000000",		-- colors: 40, 40, 40, 40
			        695 => x"00000000",		-- colors: 40, 40, 40, 40
			        696 => x"00000000",		-- colors: 40, 40, 40, 40
			        697 => x"00000000",		-- colors: 40, 40, 40, 40
			        698 => x"00000000",		-- colors: 40, 40, 40, 40
			        699 => x"00000000",		-- colors: 40, 40, 40, 40
			        700 => x"00000000",		-- colors: 40, 40, 40, 40
			        701 => x"00000000",		-- colors: 40, 40, 40, 40
			        702 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 7
			        703 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        704 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        705 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        706 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        707 => x"00000000",		-- colors: 40, 40, 40, 40
			        708 => x"00000000",		-- colors: 40, 40, 40, 40
			        709 => x"00000000",		-- colors: 40, 40, 40, 40
			        710 => x"00000000",		-- colors: 40, 40, 40, 40
			        711 => x"00000000",		-- colors: 40, 40, 40, 40
			        712 => x"00000000",		-- colors: 40, 40, 40, 40
			        713 => x"00000000",		-- colors: 40, 40, 40, 40
			        714 => x"00000000",		-- colors: 40, 40, 40, 40
			        715 => x"00000000",		-- colors: 40, 40, 40, 40
			        716 => x"00000000",		-- colors: 40, 40, 40, 40
			        717 => x"00000000",		-- colors: 40, 40, 40, 40
			        718 => x"00000000",		-- colors: 40, 40, 40, 40
			        719 => x"00000000",		-- colors: 40, 40, 40, 40
			        720 => x"00000000",		-- colors: 40, 40, 40, 40
			        721 => x"00000000",		-- colors: 40, 40, 40, 40
			        722 => x"00000000",		-- colors: 40, 40, 40, 40
			        723 => x"00000000",		-- colors: 40, 40, 40, 40
			        724 => x"00000000",		-- colors: 40, 40, 40, 40
			        725 => x"00000000",		-- colors: 40, 40, 40, 40
			        726 => x"00000000",		-- colors: 40, 40, 40, 40
			        727 => x"00000000",		-- colors: 40, 40, 40, 40
			        728 => x"00000000",		-- colors: 40, 40, 40, 40
			        729 => x"00000000",		-- colors: 40, 40, 40, 40
			        730 => x"00000000",		-- colors: 40, 40, 40, 40
			        731 => x"00000000",		-- colors: 40, 40, 40, 40
			        732 => x"00000000",		-- colors: 40, 40, 40, 40
			        733 => x"00000000",		-- colors: 40, 40, 40, 40
			        734 => x"00000000",		-- colors: 40, 40, 40, 40
			        735 => x"00000000",		-- colors: 40, 40, 40, 40
			        736 => x"00000000",		-- colors: 40, 40, 40, 40
			        737 => x"00000000",		-- colors: 40, 40, 40, 40
			        738 => x"00000000",		-- colors: 40, 40, 40, 40
			        739 => x"00000000",		-- colors: 40, 40, 40, 40
			        740 => x"00000000",		-- colors: 40, 40, 40, 40
			        741 => x"00000000",		-- colors: 40, 40, 40, 40
			        742 => x"00000000",		-- colors: 40, 40, 40, 40
			        743 => x"00000000",		-- colors: 40, 40, 40, 40
			        744 => x"00000000",		-- colors: 40, 40, 40, 40
			        745 => x"00000000",		-- colors: 40, 40, 40, 40
			        746 => x"00000000",		-- colors: 40, 40, 40, 40
			        747 => x"00000000",		-- colors: 40, 40, 40, 40
			        748 => x"00000000",		-- colors: 40, 40, 40, 40
			        749 => x"00000000",		-- colors: 40, 40, 40, 40
			        750 => x"00000000",		-- colors: 40, 40, 40, 40
			        751 => x"00000000",		-- colors: 40, 40, 40, 40
			        752 => x"00000000",		-- colors: 40, 40, 40, 40
			        753 => x"00000000",		-- colors: 40, 40, 40, 40
			        754 => x"00000000",		-- colors: 40, 40, 40, 40
			        755 => x"00000000",		-- colors: 40, 40, 40, 40
			        756 => x"00000000",		-- colors: 40, 40, 40, 40
			        757 => x"00000000",		-- colors: 40, 40, 40, 40
			        758 => x"00000000",		-- colors: 40, 40, 40, 40
			        759 => x"00000000",		-- colors: 40, 40, 40, 40
			        760 => x"00000000",		-- colors: 40, 40, 40, 40
			        761 => x"00000000",		-- colors: 40, 40, 40, 40
			        762 => x"00000000",		-- colors: 40, 40, 40, 40
			        763 => x"00000000",		-- colors: 40, 40, 40, 40
			        764 => x"00000000",		-- colors: 40, 40, 40, 40
			        765 => x"00000000",		-- colors: 40, 40, 40, 40
			        766 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 8
			        767 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        768 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        769 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        770 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        771 => x"00000000",		-- colors: 40, 40, 40, 40
			        772 => x"00000000",		-- colors: 40, 40, 40, 40
			        773 => x"00000000",		-- colors: 40, 40, 40, 40
			        774 => x"00000000",		-- colors: 40, 40, 40, 40
			        775 => x"00000000",		-- colors: 40, 40, 40, 40
			        776 => x"00000000",		-- colors: 40, 40, 40, 40
			        777 => x"00000000",		-- colors: 40, 40, 40, 40
			        778 => x"00000000",		-- colors: 40, 40, 40, 40
			        779 => x"00000000",		-- colors: 40, 40, 40, 40
			        780 => x"00000000",		-- colors: 40, 40, 40, 40
			        781 => x"00000000",		-- colors: 40, 40, 40, 40
			        782 => x"00000000",		-- colors: 40, 40, 40, 40
			        783 => x"00000000",		-- colors: 40, 40, 40, 40
			        784 => x"00000000",		-- colors: 40, 40, 40, 40
			        785 => x"00000000",		-- colors: 40, 40, 40, 40
			        786 => x"00000000",		-- colors: 40, 40, 40, 40
			        787 => x"00000000",		-- colors: 40, 40, 40, 40
			        788 => x"00000000",		-- colors: 40, 40, 40, 40
			        789 => x"00000000",		-- colors: 40, 40, 40, 40
			        790 => x"00000000",		-- colors: 40, 40, 40, 40
			        791 => x"00000000",		-- colors: 40, 40, 40, 40
			        792 => x"00000000",		-- colors: 40, 40, 40, 40
			        793 => x"00000000",		-- colors: 40, 40, 40, 40
			        794 => x"00000000",		-- colors: 40, 40, 40, 40
			        795 => x"00000000",		-- colors: 40, 40, 40, 40
			        796 => x"00000000",		-- colors: 40, 40, 40, 40
			        797 => x"00000000",		-- colors: 40, 40, 40, 40
			        798 => x"00000000",		-- colors: 40, 40, 40, 40
			        799 => x"00000000",		-- colors: 40, 40, 40, 40
			        800 => x"00000000",		-- colors: 40, 40, 40, 40
			        801 => x"00000000",		-- colors: 40, 40, 40, 40
			        802 => x"00000000",		-- colors: 40, 40, 40, 40
			        803 => x"00000000",		-- colors: 40, 40, 40, 40
			        804 => x"00000000",		-- colors: 40, 40, 40, 40
			        805 => x"00000000",		-- colors: 40, 40, 40, 40
			        806 => x"00000000",		-- colors: 40, 40, 40, 40
			        807 => x"00000000",		-- colors: 40, 40, 40, 40
			        808 => x"00000000",		-- colors: 40, 40, 40, 40
			        809 => x"00000000",		-- colors: 40, 40, 40, 40
			        810 => x"00000000",		-- colors: 40, 40, 40, 40
			        811 => x"00000000",		-- colors: 40, 40, 40, 40
			        812 => x"00000000",		-- colors: 40, 40, 40, 40
			        813 => x"00000000",		-- colors: 40, 40, 40, 40
			        814 => x"00000000",		-- colors: 40, 40, 40, 40
			        815 => x"00000000",		-- colors: 40, 40, 40, 40
			        816 => x"00000000",		-- colors: 40, 40, 40, 40
			        817 => x"00000000",		-- colors: 40, 40, 40, 40
			        818 => x"00000000",		-- colors: 40, 40, 40, 40
			        819 => x"00000000",		-- colors: 40, 40, 40, 40
			        820 => x"00000000",		-- colors: 40, 40, 40, 40
			        821 => x"00000000",		-- colors: 40, 40, 40, 40
			        822 => x"00000000",		-- colors: 40, 40, 40, 40
			        823 => x"00000000",		-- colors: 40, 40, 40, 40
			        824 => x"00000000",		-- colors: 40, 40, 40, 40
			        825 => x"00000000",		-- colors: 40, 40, 40, 40
			        826 => x"00000000",		-- colors: 40, 40, 40, 40
			        827 => x"00000000",		-- colors: 40, 40, 40, 40
			        828 => x"00000000",		-- colors: 40, 40, 40, 40
			        829 => x"00000000",		-- colors: 40, 40, 40, 40
			        830 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 9
			        831 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        832 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        833 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        834 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        835 => x"00000000",		-- colors: 40, 40, 40, 40
			        836 => x"00000000",		-- colors: 40, 40, 40, 40
			        837 => x"00000000",		-- colors: 40, 40, 40, 40
			        838 => x"00000000",		-- colors: 40, 40, 40, 40
			        839 => x"00000000",		-- colors: 40, 40, 40, 40
			        840 => x"00000000",		-- colors: 40, 40, 40, 40
			        841 => x"00000000",		-- colors: 40, 40, 40, 40
			        842 => x"00000000",		-- colors: 40, 40, 40, 40
			        843 => x"00000000",		-- colors: 40, 40, 40, 40
			        844 => x"00000000",		-- colors: 40, 40, 40, 40
			        845 => x"00000000",		-- colors: 40, 40, 40, 40
			        846 => x"00000000",		-- colors: 40, 40, 40, 40
			        847 => x"00000000",		-- colors: 40, 40, 40, 40
			        848 => x"00000000",		-- colors: 40, 40, 40, 40
			        849 => x"00000000",		-- colors: 40, 40, 40, 40
			        850 => x"00000000",		-- colors: 40, 40, 40, 40
			        851 => x"00000000",		-- colors: 40, 40, 40, 40
			        852 => x"00000000",		-- colors: 40, 40, 40, 40
			        853 => x"00000000",		-- colors: 40, 40, 40, 40
			        854 => x"00000000",		-- colors: 40, 40, 40, 40
			        855 => x"00000000",		-- colors: 40, 40, 40, 40
			        856 => x"00000000",		-- colors: 40, 40, 40, 40
			        857 => x"00000000",		-- colors: 40, 40, 40, 40
			        858 => x"00000000",		-- colors: 40, 40, 40, 40
			        859 => x"00000000",		-- colors: 40, 40, 40, 40
			        860 => x"00000000",		-- colors: 40, 40, 40, 40
			        861 => x"00000000",		-- colors: 40, 40, 40, 40
			        862 => x"00000000",		-- colors: 40, 40, 40, 40
			        863 => x"00000000",		-- colors: 40, 40, 40, 40
			        864 => x"00000000",		-- colors: 40, 40, 40, 40
			        865 => x"00000000",		-- colors: 40, 40, 40, 40
			        866 => x"00000000",		-- colors: 40, 40, 40, 40
			        867 => x"00000000",		-- colors: 40, 40, 40, 40
			        868 => x"00000000",		-- colors: 40, 40, 40, 40
			        869 => x"00000000",		-- colors: 40, 40, 40, 40
			        870 => x"00000000",		-- colors: 40, 40, 40, 40
			        871 => x"00000000",		-- colors: 40, 40, 40, 40
			        872 => x"00000000",		-- colors: 40, 40, 40, 40
			        873 => x"00000000",		-- colors: 40, 40, 40, 40
			        874 => x"00000000",		-- colors: 40, 40, 40, 40
			        875 => x"00000000",		-- colors: 40, 40, 40, 40
			        876 => x"00000000",		-- colors: 40, 40, 40, 40
			        877 => x"00000000",		-- colors: 40, 40, 40, 40
			        878 => x"00000000",		-- colors: 40, 40, 40, 40
			        879 => x"00000000",		-- colors: 40, 40, 40, 40
			        880 => x"00000000",		-- colors: 40, 40, 40, 40
			        881 => x"00000000",		-- colors: 40, 40, 40, 40
			        882 => x"00000000",		-- colors: 40, 40, 40, 40
			        883 => x"00000000",		-- colors: 40, 40, 40, 40
			        884 => x"00000000",		-- colors: 40, 40, 40, 40
			        885 => x"00000000",		-- colors: 40, 40, 40, 40
			        886 => x"00000000",		-- colors: 40, 40, 40, 40
			        887 => x"00000000",		-- colors: 40, 40, 40, 40
			        888 => x"00000000",		-- colors: 40, 40, 40, 40
			        889 => x"00000000",		-- colors: 40, 40, 40, 40
			        890 => x"00000000",		-- colors: 40, 40, 40, 40
			        891 => x"00000000",		-- colors: 40, 40, 40, 40
			        892 => x"00000000",		-- colors: 40, 40, 40, 40
			        893 => x"00000000",		-- colors: 40, 40, 40, 40
			        894 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 10
			        895 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        896 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        897 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        898 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        899 => x"00000000",		-- colors: 40, 40, 40, 40
			        900 => x"00000000",		-- colors: 40, 40, 40, 40
			        901 => x"00000000",		-- colors: 40, 40, 40, 40
			        902 => x"00000000",		-- colors: 40, 40, 40, 40
			        903 => x"00000000",		-- colors: 40, 40, 40, 40
			        904 => x"00000000",		-- colors: 40, 40, 40, 40
			        905 => x"00000000",		-- colors: 40, 40, 40, 40
			        906 => x"00000000",		-- colors: 40, 40, 40, 40
			        907 => x"00000000",		-- colors: 40, 40, 40, 40
			        908 => x"00000000",		-- colors: 40, 40, 40, 40
			        909 => x"00000000",		-- colors: 40, 40, 40, 40
			        910 => x"00000000",		-- colors: 40, 40, 40, 40
			        911 => x"00000000",		-- colors: 40, 40, 40, 40
			        912 => x"00000000",		-- colors: 40, 40, 40, 40
			        913 => x"00000000",		-- colors: 40, 40, 40, 40
			        914 => x"00000000",		-- colors: 40, 40, 40, 40
			        915 => x"00000000",		-- colors: 40, 40, 40, 40
			        916 => x"00000000",		-- colors: 40, 40, 40, 40
			        917 => x"00000000",		-- colors: 40, 40, 40, 40
			        918 => x"00000000",		-- colors: 40, 40, 40, 40
			        919 => x"00000000",		-- colors: 40, 40, 40, 40
			        920 => x"00000000",		-- colors: 40, 40, 40, 40
			        921 => x"00000000",		-- colors: 40, 40, 40, 40
			        922 => x"00000000",		-- colors: 40, 40, 40, 40
			        923 => x"00000000",		-- colors: 40, 40, 40, 40
			        924 => x"00000000",		-- colors: 40, 40, 40, 40
			        925 => x"00000000",		-- colors: 40, 40, 40, 40
			        926 => x"00000000",		-- colors: 40, 40, 40, 40
			        927 => x"00000000",		-- colors: 40, 40, 40, 40
			        928 => x"00000000",		-- colors: 40, 40, 40, 40
			        929 => x"00000000",		-- colors: 40, 40, 40, 40
			        930 => x"00000000",		-- colors: 40, 40, 40, 40
			        931 => x"00000000",		-- colors: 40, 40, 40, 40
			        932 => x"00000000",		-- colors: 40, 40, 40, 40
			        933 => x"00000000",		-- colors: 40, 40, 40, 40
			        934 => x"00000000",		-- colors: 40, 40, 40, 40
			        935 => x"00000000",		-- colors: 40, 40, 40, 40
			        936 => x"00000000",		-- colors: 40, 40, 40, 40
			        937 => x"00000000",		-- colors: 40, 40, 40, 40
			        938 => x"00000000",		-- colors: 40, 40, 40, 40
			        939 => x"00000000",		-- colors: 40, 40, 40, 40
			        940 => x"00000000",		-- colors: 40, 40, 40, 40
			        941 => x"00000000",		-- colors: 40, 40, 40, 40
			        942 => x"00000000",		-- colors: 40, 40, 40, 40
			        943 => x"00000000",		-- colors: 40, 40, 40, 40
			        944 => x"00000000",		-- colors: 40, 40, 40, 40
			        945 => x"00000000",		-- colors: 40, 40, 40, 40
			        946 => x"00000000",		-- colors: 40, 40, 40, 40
			        947 => x"00000000",		-- colors: 40, 40, 40, 40
			        948 => x"00000000",		-- colors: 40, 40, 40, 40
			        949 => x"00000000",		-- colors: 40, 40, 40, 40
			        950 => x"00000000",		-- colors: 40, 40, 40, 40
			        951 => x"00000000",		-- colors: 40, 40, 40, 40
			        952 => x"00000000",		-- colors: 40, 40, 40, 40
			        953 => x"00000000",		-- colors: 40, 40, 40, 40
			        954 => x"00000000",		-- colors: 40, 40, 40, 40
			        955 => x"00000000",		-- colors: 40, 40, 40, 40
			        956 => x"00000000",		-- colors: 40, 40, 40, 40
			        957 => x"00000000",		-- colors: 40, 40, 40, 40
			        958 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 11
			        959 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        960 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        961 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        962 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        963 => x"00000000",		-- colors: 40, 40, 40, 40
			        964 => x"00000000",		-- colors: 40, 40, 40, 40
			        965 => x"00000000",		-- colors: 40, 40, 40, 40
			        966 => x"00000000",		-- colors: 40, 40, 40, 40
			        967 => x"00000000",		-- colors: 40, 40, 40, 40
			        968 => x"00000000",		-- colors: 40, 40, 40, 40
			        969 => x"00000000",		-- colors: 40, 40, 40, 40
			        970 => x"00000000",		-- colors: 40, 40, 40, 40
			        971 => x"00000000",		-- colors: 40, 40, 40, 40
			        972 => x"00000000",		-- colors: 40, 40, 40, 40
			        973 => x"00000000",		-- colors: 40, 40, 40, 40
			        974 => x"00000000",		-- colors: 40, 40, 40, 40
			        975 => x"00000000",		-- colors: 40, 40, 40, 40
			        976 => x"00000000",		-- colors: 40, 40, 40, 40
			        977 => x"00000000",		-- colors: 40, 40, 40, 40
			        978 => x"00000000",		-- colors: 40, 40, 40, 40
			        979 => x"00000000",		-- colors: 40, 40, 40, 40
			        980 => x"00000000",		-- colors: 40, 40, 40, 40
			        981 => x"00000000",		-- colors: 40, 40, 40, 40
			        982 => x"00000000",		-- colors: 40, 40, 40, 40
			        983 => x"00000000",		-- colors: 40, 40, 40, 40
			        984 => x"00000000",		-- colors: 40, 40, 40, 40
			        985 => x"00000000",		-- colors: 40, 40, 40, 40
			        986 => x"00000000",		-- colors: 40, 40, 40, 40
			        987 => x"00000000",		-- colors: 40, 40, 40, 40
			        988 => x"00000000",		-- colors: 40, 40, 40, 40
			        989 => x"00000000",		-- colors: 40, 40, 40, 40
			        990 => x"00000000",		-- colors: 40, 40, 40, 40
			        991 => x"00000000",		-- colors: 40, 40, 40, 40
			        992 => x"00000000",		-- colors: 40, 40, 40, 40
			        993 => x"00000000",		-- colors: 40, 40, 40, 40
			        994 => x"00000000",		-- colors: 40, 40, 40, 40
			        995 => x"00000000",		-- colors: 40, 40, 40, 40
			        996 => x"00000000",		-- colors: 40, 40, 40, 40
			        997 => x"00000000",		-- colors: 40, 40, 40, 40
			        998 => x"00000000",		-- colors: 40, 40, 40, 40
			        999 => x"00000000",		-- colors: 40, 40, 40, 40
			        1000 => x"00000000",		-- colors: 40, 40, 40, 40
			        1001 => x"00000000",		-- colors: 40, 40, 40, 40
			        1002 => x"00000000",		-- colors: 40, 40, 40, 40
			        1003 => x"00000000",		-- colors: 40, 40, 40, 40
			        1004 => x"00000000",		-- colors: 40, 40, 40, 40
			        1005 => x"00000000",		-- colors: 40, 40, 40, 40
			        1006 => x"00000000",		-- colors: 40, 40, 40, 40
			        1007 => x"00000000",		-- colors: 40, 40, 40, 40
			        1008 => x"00000000",		-- colors: 40, 40, 40, 40
			        1009 => x"00000000",		-- colors: 40, 40, 40, 40
			        1010 => x"00000000",		-- colors: 40, 40, 40, 40
			        1011 => x"00000000",		-- colors: 40, 40, 40, 40
			        1012 => x"00000000",		-- colors: 40, 40, 40, 40
			        1013 => x"00000000",		-- colors: 40, 40, 40, 40
			        1014 => x"00000000",		-- colors: 40, 40, 40, 40
			        1015 => x"00000000",		-- colors: 40, 40, 40, 40
			        1016 => x"00000000",		-- colors: 40, 40, 40, 40
			        1017 => x"00000000",		-- colors: 40, 40, 40, 40
			        1018 => x"00000000",		-- colors: 40, 40, 40, 40
			        1019 => x"00000000",		-- colors: 40, 40, 40, 40
			        1020 => x"00000000",		-- colors: 40, 40, 40, 40
			        1021 => x"00000000",		-- colors: 40, 40, 40, 40
			        1022 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 12
			        1023 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        1024 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        1025 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        1026 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        1027 => x"00000000",		-- colors: 40, 40, 40, 40
			        1028 => x"00000000",		-- colors: 40, 40, 40, 40
			        1029 => x"00000000",		-- colors: 40, 40, 40, 40
			        1030 => x"00000000",		-- colors: 40, 40, 40, 40
			        1031 => x"00000000",		-- colors: 40, 40, 40, 40
			        1032 => x"00000000",		-- colors: 40, 40, 40, 40
			        1033 => x"00000000",		-- colors: 40, 40, 40, 40
			        1034 => x"00000000",		-- colors: 40, 40, 40, 40
			        1035 => x"00000000",		-- colors: 40, 40, 40, 40
			        1036 => x"00000000",		-- colors: 40, 40, 40, 40
			        1037 => x"00000000",		-- colors: 40, 40, 40, 40
			        1038 => x"00000000",		-- colors: 40, 40, 40, 40
			        1039 => x"00000000",		-- colors: 40, 40, 40, 40
			        1040 => x"00000000",		-- colors: 40, 40, 40, 40
			        1041 => x"00000000",		-- colors: 40, 40, 40, 40
			        1042 => x"00000000",		-- colors: 40, 40, 40, 40
			        1043 => x"00000000",		-- colors: 40, 40, 40, 40
			        1044 => x"00000000",		-- colors: 40, 40, 40, 40
			        1045 => x"00000000",		-- colors: 40, 40, 40, 40
			        1046 => x"00000000",		-- colors: 40, 40, 40, 40
			        1047 => x"00000000",		-- colors: 40, 40, 40, 40
			        1048 => x"00000000",		-- colors: 40, 40, 40, 40
			        1049 => x"00000000",		-- colors: 40, 40, 40, 40
			        1050 => x"00000000",		-- colors: 40, 40, 40, 40
			        1051 => x"00000000",		-- colors: 40, 40, 40, 40
			        1052 => x"00000000",		-- colors: 40, 40, 40, 40
			        1053 => x"00000000",		-- colors: 40, 40, 40, 40
			        1054 => x"00000000",		-- colors: 40, 40, 40, 40
			        1055 => x"00000000",		-- colors: 40, 40, 40, 40
			        1056 => x"00000000",		-- colors: 40, 40, 40, 40
			        1057 => x"00000000",		-- colors: 40, 40, 40, 40
			        1058 => x"00000000",		-- colors: 40, 40, 40, 40
			        1059 => x"00000000",		-- colors: 40, 40, 40, 40
			        1060 => x"00000000",		-- colors: 40, 40, 40, 40
			        1061 => x"00000000",		-- colors: 40, 40, 40, 40
			        1062 => x"00000000",		-- colors: 40, 40, 40, 40
			        1063 => x"00000000",		-- colors: 40, 40, 40, 40
			        1064 => x"00000000",		-- colors: 40, 40, 40, 40
			        1065 => x"00000000",		-- colors: 40, 40, 40, 40
			        1066 => x"00000000",		-- colors: 40, 40, 40, 40
			        1067 => x"00000000",		-- colors: 40, 40, 40, 40
			        1068 => x"00000000",		-- colors: 40, 40, 40, 40
			        1069 => x"00000000",		-- colors: 40, 40, 40, 40
			        1070 => x"00000000",		-- colors: 40, 40, 40, 40
			        1071 => x"00000000",		-- colors: 40, 40, 40, 40
			        1072 => x"00000000",		-- colors: 40, 40, 40, 40
			        1073 => x"00000000",		-- colors: 40, 40, 40, 40
			        1074 => x"00000000",		-- colors: 40, 40, 40, 40
			        1075 => x"00000000",		-- colors: 40, 40, 40, 40
			        1076 => x"00000000",		-- colors: 40, 40, 40, 40
			        1077 => x"00000000",		-- colors: 40, 40, 40, 40
			        1078 => x"00000000",		-- colors: 40, 40, 40, 40
			        1079 => x"00000000",		-- colors: 40, 40, 40, 40
			        1080 => x"00000000",		-- colors: 40, 40, 40, 40
			        1081 => x"00000000",		-- colors: 40, 40, 40, 40
			        1082 => x"00000000",		-- colors: 40, 40, 40, 40
			        1083 => x"00000000",		-- colors: 40, 40, 40, 40
			        1084 => x"00000000",		-- colors: 40, 40, 40, 40
			        1085 => x"00000000",		-- colors: 40, 40, 40, 40
			        1086 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 13
			        1087 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        1088 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        1089 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        1090 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        1091 => x"00000000",		-- colors: 40, 40, 40, 40
			        1092 => x"00000000",		-- colors: 40, 40, 40, 40
			        1093 => x"00000000",		-- colors: 40, 40, 40, 40
			        1094 => x"00000000",		-- colors: 40, 40, 40, 40
			        1095 => x"00000000",		-- colors: 40, 40, 40, 40
			        1096 => x"00000000",		-- colors: 40, 40, 40, 40
			        1097 => x"00000000",		-- colors: 40, 40, 40, 40
			        1098 => x"00000000",		-- colors: 40, 40, 40, 40
			        1099 => x"00000000",		-- colors: 40, 40, 40, 40
			        1100 => x"00000000",		-- colors: 40, 40, 40, 40
			        1101 => x"00000000",		-- colors: 40, 40, 40, 40
			        1102 => x"00000000",		-- colors: 40, 40, 40, 40
			        1103 => x"00000000",		-- colors: 40, 40, 40, 40
			        1104 => x"00000000",		-- colors: 40, 40, 40, 40
			        1105 => x"00000000",		-- colors: 40, 40, 40, 40
			        1106 => x"00000000",		-- colors: 40, 40, 40, 40
			        1107 => x"00000000",		-- colors: 40, 40, 40, 40
			        1108 => x"00000000",		-- colors: 40, 40, 40, 40
			        1109 => x"00000000",		-- colors: 40, 40, 40, 40
			        1110 => x"00000000",		-- colors: 40, 40, 40, 40
			        1111 => x"00000000",		-- colors: 40, 40, 40, 40
			        1112 => x"00000000",		-- colors: 40, 40, 40, 40
			        1113 => x"00000000",		-- colors: 40, 40, 40, 40
			        1114 => x"00000000",		-- colors: 40, 40, 40, 40
			        1115 => x"00000000",		-- colors: 40, 40, 40, 40
			        1116 => x"00000000",		-- colors: 40, 40, 40, 40
			        1117 => x"00000000",		-- colors: 40, 40, 40, 40
			        1118 => x"00000000",		-- colors: 40, 40, 40, 40
			        1119 => x"00000000",		-- colors: 40, 40, 40, 40
			        1120 => x"00000000",		-- colors: 40, 40, 40, 40
			        1121 => x"00000000",		-- colors: 40, 40, 40, 40
			        1122 => x"00000000",		-- colors: 40, 40, 40, 40
			        1123 => x"00000000",		-- colors: 40, 40, 40, 40
			        1124 => x"00000000",		-- colors: 40, 40, 40, 40
			        1125 => x"00000000",		-- colors: 40, 40, 40, 40
			        1126 => x"00000000",		-- colors: 40, 40, 40, 40
			        1127 => x"00000000",		-- colors: 40, 40, 40, 40
			        1128 => x"00000000",		-- colors: 40, 40, 40, 40
			        1129 => x"00000000",		-- colors: 40, 40, 40, 40
			        1130 => x"00000000",		-- colors: 40, 40, 40, 40
			        1131 => x"00000000",		-- colors: 40, 40, 40, 40
			        1132 => x"00000000",		-- colors: 40, 40, 40, 40
			        1133 => x"00000000",		-- colors: 40, 40, 40, 40
			        1134 => x"00000000",		-- colors: 40, 40, 40, 40
			        1135 => x"00000000",		-- colors: 40, 40, 40, 40
			        1136 => x"00000000",		-- colors: 40, 40, 40, 40
			        1137 => x"00000000",		-- colors: 40, 40, 40, 40
			        1138 => x"00000000",		-- colors: 40, 40, 40, 40
			        1139 => x"00000000",		-- colors: 40, 40, 40, 40
			        1140 => x"00000000",		-- colors: 40, 40, 40, 40
			        1141 => x"00000000",		-- colors: 40, 40, 40, 40
			        1142 => x"00000000",		-- colors: 40, 40, 40, 40
			        1143 => x"00000000",		-- colors: 40, 40, 40, 40
			        1144 => x"00000000",		-- colors: 40, 40, 40, 40
			        1145 => x"00000000",		-- colors: 40, 40, 40, 40
			        1146 => x"00000000",		-- colors: 40, 40, 40, 40
			        1147 => x"00000000",		-- colors: 40, 40, 40, 40
			        1148 => x"00000000",		-- colors: 40, 40, 40, 40
			        1149 => x"00000000",		-- colors: 40, 40, 40, 40
			        1150 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 14
			        1151 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        1152 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        1153 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        1154 => x"2C2C2C2C",		-- colors: 44, 44, 44, 44
			        1155 => x"00000000",		-- colors: 40, 40, 40, 40
			        1156 => x"00000000",		-- colors: 40, 40, 40, 40
			        1157 => x"00000000",		-- colors: 40, 40, 40, 40
			        1158 => x"00000000",		-- colors: 40, 40, 40, 40
			        1159 => x"00000000",		-- colors: 40, 40, 40, 40
			        1160 => x"00000000",		-- colors: 40, 40, 40, 40
			        1161 => x"00000000",		-- colors: 40, 40, 40, 40
			        1162 => x"00000000",		-- colors: 40, 40, 40, 40
			        1163 => x"00000000",		-- colors: 40, 40, 40, 40
			        1164 => x"00000000",		-- colors: 40, 40, 40, 40
			        1165 => x"00000000",		-- colors: 40, 40, 40, 40
			        1166 => x"00000000",		-- colors: 40, 40, 40, 40
			        1167 => x"00000000",		-- colors: 40, 40, 40, 40
			        1168 => x"00000000",		-- colors: 40, 40, 40, 40
			        1169 => x"00000000",		-- colors: 40, 40, 40, 40
			        1170 => x"00000000",		-- colors: 40, 40, 40, 40
			        1171 => x"00000000",		-- colors: 40, 40, 40, 40
			        1172 => x"00000000",		-- colors: 40, 40, 40, 40
			        1173 => x"00000000",		-- colors: 40, 40, 40, 40
			        1174 => x"00000000",		-- colors: 40, 40, 40, 40
			        1175 => x"00000000",		-- colors: 40, 40, 40, 40
			        1176 => x"00000000",		-- colors: 40, 40, 40, 40
			        1177 => x"00000000",		-- colors: 40, 40, 40, 40
			        1178 => x"00000000",		-- colors: 40, 40, 40, 40
			        1179 => x"00000000",		-- colors: 40, 40, 40, 40
			        1180 => x"00000000",		-- colors: 40, 40, 40, 40
			        1181 => x"00000000",		-- colors: 40, 40, 40, 40
			        1182 => x"00000000",		-- colors: 40, 40, 40, 40
			        1183 => x"00000000",		-- colors: 40, 40, 40, 40
			        1184 => x"00000000",		-- colors: 40, 40, 40, 40
			        1185 => x"00000000",		-- colors: 40, 40, 40, 40
			        1186 => x"00000000",		-- colors: 40, 40, 40, 40
			        1187 => x"00000000",		-- colors: 40, 40, 40, 40
			        1188 => x"00000000",		-- colors: 40, 40, 40, 40
			        1189 => x"00000000",		-- colors: 40, 40, 40, 40
			        1190 => x"00000000",		-- colors: 40, 40, 40, 40
			        1191 => x"00000000",		-- colors: 40, 40, 40, 40
			        1192 => x"00000000",		-- colors: 40, 40, 40, 40
			        1193 => x"00000000",		-- colors: 40, 40, 40, 40
			        1194 => x"00000000",		-- colors: 40, 40, 40, 40
			        1195 => x"00000000",		-- colors: 40, 40, 40, 40
			        1196 => x"00000000",		-- colors: 40, 40, 40, 40
			        1197 => x"00000000",		-- colors: 40, 40, 40, 40
			        1198 => x"00000000",		-- colors: 40, 40, 40, 40
			        1199 => x"00000000",		-- colors: 40, 40, 40, 40
			        1200 => x"00000000",		-- colors: 40, 40, 40, 40
			        1201 => x"00000000",		-- colors: 40, 40, 40, 40
			        1202 => x"00000000",		-- colors: 40, 40, 40, 40
			        1203 => x"00000000",		-- colors: 40, 40, 40, 40
			        1204 => x"00000000",		-- colors: 40, 40, 40, 40
			        1205 => x"00000000",		-- colors: 40, 40, 40, 40
			        1206 => x"00000000",		-- colors: 40, 40, 40, 40
			        1207 => x"00000000",		-- colors: 40, 40, 40, 40
			        1208 => x"00000000",		-- colors: 40, 40, 40, 40
			        1209 => x"00000000",		-- colors: 40, 40, 40, 40
			        1210 => x"00000000",		-- colors: 40, 40, 40, 40
			        1211 => x"00000000",		-- colors: 40, 40, 40, 40
			        1212 => x"00000000",		-- colors: 40, 40, 40, 40
			        1213 => x"00000000",		-- colors: 40, 40, 40, 40
			        1214 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 15
			        1215 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
			        1216 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
			        1217 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
			        1218 => x"2D2D2D2D",		-- colors: 45, 45, 45, 45
			        1219 => x"00000000",		-- colors: 40, 40, 40, 40
			        1220 => x"00000000",		-- colors: 40, 40, 40, 40
			        1221 => x"00000000",		-- colors: 40, 40, 40, 40
			        1222 => x"00000000",		-- colors: 40, 40, 40, 40
			        1223 => x"00000000",		-- colors: 40, 40, 40, 40
			        1224 => x"00000000",		-- colors: 40, 40, 40, 40
			        1225 => x"00000000",		-- colors: 40, 40, 40, 40
			        1226 => x"00000000",		-- colors: 40, 40, 40, 40
			        1227 => x"00000000",		-- colors: 40, 40, 40, 40
			        1228 => x"00000000",		-- colors: 40, 40, 40, 40
			        1229 => x"00000000",		-- colors: 40, 40, 40, 40
			        1230 => x"00000000",		-- colors: 40, 40, 40, 40
			        1231 => x"00000000",		-- colors: 40, 40, 40, 40
			        1232 => x"00000000",		-- colors: 40, 40, 40, 40
			        1233 => x"00000000",		-- colors: 40, 40, 40, 40
			        1234 => x"00000000",		-- colors: 40, 40, 40, 40
			        1235 => x"00000000",		-- colors: 40, 40, 40, 40
			        1236 => x"00000000",		-- colors: 40, 40, 40, 40
			        1237 => x"00000000",		-- colors: 40, 40, 40, 40
			        1238 => x"00000000",		-- colors: 40, 40, 40, 40
			        1239 => x"00000000",		-- colors: 40, 40, 40, 40
			        1240 => x"00000000",		-- colors: 40, 40, 40, 40
			        1241 => x"00000000",		-- colors: 40, 40, 40, 40
			        1242 => x"00000000",		-- colors: 40, 40, 40, 40
			        1243 => x"00000000",		-- colors: 40, 40, 40, 40
			        1244 => x"00000000",		-- colors: 40, 40, 40, 40
			        1245 => x"00000000",		-- colors: 40, 40, 40, 40
			        1246 => x"00000000",		-- colors: 40, 40, 40, 40
			        1247 => x"00000000",		-- colors: 40, 40, 40, 40
			        1248 => x"00000000",		-- colors: 40, 40, 40, 40
			        1249 => x"00000000",		-- colors: 40, 40, 40, 40
			        1250 => x"00000000",		-- colors: 40, 40, 40, 40
			        1251 => x"00000000",		-- colors: 40, 40, 40, 40
			        1252 => x"00000000",		-- colors: 40, 40, 40, 40
			        1253 => x"00000000",		-- colors: 40, 40, 40, 40
			        1254 => x"00000000",		-- colors: 40, 40, 40, 40
			        1255 => x"00000000",		-- colors: 40, 40, 40, 40
			        1256 => x"00000000",		-- colors: 40, 40, 40, 40
			        1257 => x"00000000",		-- colors: 40, 40, 40, 40
			        1258 => x"00000000",		-- colors: 40, 40, 40, 40
			        1259 => x"00000000",		-- colors: 40, 40, 40, 40
			        1260 => x"00000000",		-- colors: 40, 40, 40, 40
			        1261 => x"00000000",		-- colors: 40, 40, 40, 40
			        1262 => x"00000000",		-- colors: 40, 40, 40, 40
			        1263 => x"00000000",		-- colors: 40, 40, 40, 40
			        1264 => x"00000000",		-- colors: 40, 40, 40, 40
			        1265 => x"00000000",		-- colors: 40, 40, 40, 40
			        1266 => x"00000000",		-- colors: 40, 40, 40, 40
			        1267 => x"00000000",		-- colors: 40, 40, 40, 40
			        1268 => x"00000000",		-- colors: 40, 40, 40, 40
			        1269 => x"00000000",		-- colors: 40, 40, 40, 40
			        1270 => x"00000000",		-- colors: 40, 40, 40, 40
			        1271 => x"00000000",		-- colors: 40, 40, 40, 40
			        1272 => x"00000000",		-- colors: 40, 40, 40, 40
			        1273 => x"00000000",		-- colors: 40, 40, 40, 40
			        1274 => x"00000000",		-- colors: 40, 40, 40, 40
			        1275 => x"00000000",		-- colors: 40, 40, 40, 40
			        1276 => x"00000000",		-- colors: 40, 40, 40, 40
			        1277 => x"00000000",		-- colors: 40, 40, 40, 40
			        1278 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 16
			        1279 => x"00000000",		-- colors: 40, 40, 40, 40
			        1280 => x"00000000",		-- colors: 40, 40, 40, 40
			        1281 => x"00000000",		-- colors: 40, 40, 40, 40
			        1282 => x"00000000",		-- colors: 40, 40, 40, 40
			        1283 => x"00000000",		-- colors: 40, 40, 40, 40
			        1284 => x"00000000",		-- colors: 40, 40, 40, 40
			        1285 => x"00000000",		-- colors: 40, 40, 40, 40
			        1286 => x"00000000",		-- colors: 40, 40, 40, 40
			        1287 => x"00000000",		-- colors: 40, 40, 40, 40
			        1288 => x"00000000",		-- colors: 40, 40, 40, 40
			        1289 => x"00000000",		-- colors: 40, 40, 40, 40
			        1290 => x"00000000",		-- colors: 40, 40, 40, 40
			        1291 => x"00000000",		-- colors: 40, 40, 40, 40
			        1292 => x"00000000",		-- colors: 40, 40, 40, 40
			        1293 => x"00000000",		-- colors: 40, 40, 40, 40
			        1294 => x"00000000",		-- colors: 40, 40, 40, 40
			        1295 => x"00000000",		-- colors: 40, 40, 40, 40
			        1296 => x"00000000",		-- colors: 40, 40, 40, 40
			        1297 => x"00000000",		-- colors: 40, 40, 40, 40
			        1298 => x"00000000",		-- colors: 40, 40, 40, 40
			        1299 => x"00000000",		-- colors: 40, 40, 40, 40
			        1300 => x"00000000",		-- colors: 40, 40, 40, 40
			        1301 => x"00000000",		-- colors: 40, 40, 40, 40
			        1302 => x"00000000",		-- colors: 40, 40, 40, 40
			        1303 => x"00000000",		-- colors: 40, 40, 40, 40
			        1304 => x"00000000",		-- colors: 40, 40, 40, 40
			        1305 => x"00000000",		-- colors: 40, 40, 40, 40
			        1306 => x"00000000",		-- colors: 40, 40, 40, 40
			        1307 => x"00000000",		-- colors: 40, 40, 40, 40
			        1308 => x"00000000",		-- colors: 40, 40, 40, 40
			        1309 => x"00000000",		-- colors: 40, 40, 40, 40
			        1310 => x"00000000",		-- colors: 40, 40, 40, 40
			        1311 => x"00000000",		-- colors: 40, 40, 40, 40
			        1312 => x"00000000",		-- colors: 40, 40, 40, 40
			        1313 => x"00000000",		-- colors: 40, 40, 40, 40
			        1314 => x"00000000",		-- colors: 40, 40, 40, 40
			        1315 => x"00000000",		-- colors: 40, 40, 40, 40
			        1316 => x"00000000",		-- colors: 40, 40, 40, 40
			        1317 => x"00000000",		-- colors: 40, 40, 40, 40
			        1318 => x"00000000",		-- colors: 40, 40, 40, 40
			        1319 => x"00000000",		-- colors: 40, 40, 40, 40
			        1320 => x"00000000",		-- colors: 40, 40, 40, 40
			        1321 => x"00000000",		-- colors: 40, 40, 40, 40
			        1322 => x"00000000",		-- colors: 40, 40, 40, 40
			        1323 => x"00000000",		-- colors: 40, 40, 40, 40
			        1324 => x"00000000",		-- colors: 40, 40, 40, 40
			        1325 => x"00000000",		-- colors: 40, 40, 40, 40
			        1326 => x"00000000",		-- colors: 40, 40, 40, 40
			        1327 => x"00000000",		-- colors: 40, 40, 40, 40
			        1328 => x"00000000",		-- colors: 40, 40, 40, 40
			        1329 => x"00000000",		-- colors: 40, 40, 40, 40
			        1330 => x"00000000",		-- colors: 40, 40, 40, 40
			        1331 => x"00000000",		-- colors: 40, 40, 40, 40
			        1332 => x"00000000",		-- colors: 40, 40, 40, 40
			        1333 => x"00000000",		-- colors: 40, 40, 40, 40
			        1334 => x"00000000",		-- colors: 40, 40, 40, 40
			        1335 => x"00000000",		-- colors: 40, 40, 40, 40
			        1336 => x"00000000",		-- colors: 40, 40, 40, 40
			        1337 => x"00000000",		-- colors: 40, 40, 40, 40
			        1338 => x"00000000",		-- colors: 40, 40, 40, 40
			        1339 => x"36363636",		-- colors: 54, 54, 54, 54
			        1340 => x"36363636",		-- colors: 54, 54, 54, 54
			        1341 => x"36363636",		-- colors: 54, 54, 54, 54
			        1342 => x"36363636",		-- colors: 54, 54, 54, 54

			                --  sprite 17
			        1343 => x"00000000",		-- colors: 40, 40, 40, 40
			        1344 => x"00000000",		-- colors: 40, 40, 40, 40
			        1345 => x"00000000",		-- colors: 40, 40, 40, 40
			        1346 => x"00000000",		-- colors: 40, 40, 40, 40
			        1347 => x"3A3A3A3A",		-- colors: 58, 58, 58, 58
			        1348 => x"3A3A3A3A",		-- colors: 58, 58, 58, 58
			        1349 => x"3A3A3A3A",		-- colors: 58, 58, 58, 58
			        1350 => x"3A3A3A3A",		-- colors: 58, 58, 58, 58
			        1351 => x"3B3B3B3B",		-- colors: 59, 59, 59, 59
			        1352 => x"3B3B3B3B",		-- colors: 59, 59, 59, 59
			        1353 => x"3B3B3B3B",		-- colors: 59, 59, 59, 59
			        1354 => x"3B3B3B3B",		-- colors: 59, 59, 59, 59
			        1355 => x"39393939",		-- colors: 57, 57, 57, 57
			        1356 => x"39393939",		-- colors: 57, 57, 57, 57
			        1357 => x"39393939",		-- colors: 57, 57, 57, 57
			        1358 => x"39393939",		-- colors: 57, 57, 57, 57
			        1359 => x"39393939",		-- colors: 57, 57, 57, 57
			        1360 => x"39393939",		-- colors: 57, 57, 57, 57
			        1361 => x"39393939",		-- colors: 57, 57, 57, 57
			        1362 => x"39393939",		-- colors: 57, 57, 57, 57
			        1363 => x"39393939",		-- colors: 57, 57, 57, 57
			        1364 => x"39393939",		-- colors: 57, 57, 57, 57
			        1365 => x"39393939",		-- colors: 57, 57, 57, 57
			        1366 => x"39393939",		-- colors: 57, 57, 57, 57
			        1367 => x"39393939",		-- colors: 57, 57, 57, 57
			        1368 => x"39393939",		-- colors: 57, 57, 57, 57
			        1369 => x"39393939",		-- colors: 57, 57, 57, 57
			        1370 => x"39393939",		-- colors: 57, 57, 57, 57
			        1371 => x"39393939",		-- colors: 57, 57, 57, 57
			        1372 => x"39393939",		-- colors: 57, 57, 57, 57
			        1373 => x"39393939",		-- colors: 57, 57, 57, 57
			        1374 => x"39393939",		-- colors: 57, 57, 57, 57
			        1375 => x"39393939",		-- colors: 57, 57, 57, 57
			        1376 => x"39393939",		-- colors: 57, 57, 57, 57
			        1377 => x"39393939",		-- colors: 57, 57, 57, 57
			        1378 => x"39393939",		-- colors: 57, 57, 57, 57
			        1379 => x"39393939",		-- colors: 57, 57, 57, 57
			        1380 => x"39393939",		-- colors: 57, 57, 57, 57
			        1381 => x"39393939",		-- colors: 57, 57, 57, 57
			        1382 => x"39393939",		-- colors: 57, 57, 57, 57
			        1383 => x"39393939",		-- colors: 57, 57, 57, 57
			        1384 => x"39393939",		-- colors: 57, 57, 57, 57
			        1385 => x"39393939",		-- colors: 57, 57, 57, 57
			        1386 => x"39393939",		-- colors: 57, 57, 57, 57
			        1387 => x"39393939",		-- colors: 57, 57, 57, 57
			        1388 => x"39393939",		-- colors: 57, 57, 57, 57
			        1389 => x"39393939",		-- colors: 57, 57, 57, 57
			        1390 => x"39393939",		-- colors: 57, 57, 57, 57
			        1391 => x"39393939",		-- colors: 57, 57, 57, 57
			        1392 => x"39393939",		-- colors: 57, 57, 57, 57
			        1393 => x"39393939",		-- colors: 57, 57, 57, 57
			        1394 => x"39393939",		-- colors: 57, 57, 57, 57
			        1395 => x"39393939",		-- colors: 57, 57, 57, 57
			        1396 => x"39393939",		-- colors: 57, 57, 57, 57
			        1397 => x"39393939",		-- colors: 57, 57, 57, 57
			        1398 => x"39393939",		-- colors: 57, 57, 57, 57
			        1399 => x"39393939",		-- colors: 57, 57, 57, 57
			        1400 => x"39393939",		-- colors: 57, 57, 57, 57
			        1401 => x"39393939",		-- colors: 57, 57, 57, 57
			        1402 => x"39393939",		-- colors: 57, 57, 57, 57
			        1403 => x"3B3B3B3B",		-- colors: 59, 59, 59, 59
			        1404 => x"3B3B3B3B",		-- colors: 59, 59, 59, 59
			        1405 => x"3B3B3B3B",		-- colors: 59, 59, 59, 59
			        1406 => x"3B3B3B3B",		-- colors: 59, 59, 59, 59

			                --  sprite 18
			        1407 => x"00000000",		-- colors: 40, 40, 40, 40
			        1408 => x"00000000",		-- colors: 40, 40, 40, 40
			        1409 => x"00000000",		-- colors: 40, 40, 40, 40
			        1410 => x"00000000",		-- colors: 40, 40, 40, 40
			        1411 => x"00000000",		-- colors: 40, 40, 40, 40
			        1412 => x"00000000",		-- colors: 40, 40, 40, 40
			        1413 => x"00000000",		-- colors: 40, 40, 40, 40
			        1414 => x"00000000",		-- colors: 40, 40, 40, 40
			        1415 => x"00000000",		-- colors: 40, 40, 40, 40
			        1416 => x"00000000",		-- colors: 40, 40, 40, 40
			        1417 => x"00000000",		-- colors: 40, 40, 40, 40
			        1418 => x"00000000",		-- colors: 40, 40, 40, 40
			        1419 => x"00000000",		-- colors: 40, 40, 40, 40
			        1420 => x"00000000",		-- colors: 40, 40, 40, 40
			        1421 => x"00000000",		-- colors: 40, 40, 40, 40
			        1422 => x"00000000",		-- colors: 40, 40, 40, 40
			        1423 => x"00000000",		-- colors: 40, 40, 40, 40
			        1424 => x"00000000",		-- colors: 40, 40, 40, 40
			        1425 => x"00000000",		-- colors: 40, 40, 40, 40
			        1426 => x"00000000",		-- colors: 40, 40, 40, 40
			        1427 => x"00000000",		-- colors: 40, 40, 40, 40
			        1428 => x"00000000",		-- colors: 40, 40, 40, 40
			        1429 => x"00000000",		-- colors: 40, 40, 40, 40
			        1430 => x"00000000",		-- colors: 40, 40, 40, 40
			        1431 => x"00000000",		-- colors: 40, 40, 40, 40
			        1432 => x"00000000",		-- colors: 40, 40, 40, 40
			        1433 => x"00000000",		-- colors: 40, 40, 40, 40
			        1434 => x"00000000",		-- colors: 40, 40, 40, 40
			        1435 => x"00000000",		-- colors: 40, 40, 40, 40
			        1436 => x"00000000",		-- colors: 40, 40, 40, 40
			        1437 => x"00000000",		-- colors: 40, 40, 40, 40
			        1438 => x"00000000",		-- colors: 40, 40, 40, 40
			        1439 => x"00000000",		-- colors: 40, 40, 40, 40
			        1440 => x"00000000",		-- colors: 40, 40, 40, 40
			        1441 => x"00000000",		-- colors: 40, 40, 40, 40
			        1442 => x"00000000",		-- colors: 40, 40, 40, 40
			        1443 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1444 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1445 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1446 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1447 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1448 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1449 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1450 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1451 => x"00000000",		-- colors: 40, 40, 40, 40
			        1452 => x"00000000",		-- colors: 40, 40, 40, 40
			        1453 => x"00000000",		-- colors: 40, 40, 40, 40
			        1454 => x"00000000",		-- colors: 40, 40, 40, 40
			        1455 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1456 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1457 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1458 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1459 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1460 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1461 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1462 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1463 => x"00000000",		-- colors: 40, 40, 40, 40
			        1464 => x"00000000",		-- colors: 40, 40, 40, 40
			        1465 => x"00000000",		-- colors: 40, 40, 40, 40
			        1466 => x"00000000",		-- colors: 40, 40, 40, 40
			        1467 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1468 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1469 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1470 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60

			                --  sprite 19
			        1471 => x"00000000",		-- colors: 40, 40, 40, 40
			        1472 => x"00000000",		-- colors: 40, 40, 40, 40
			        1473 => x"00000000",		-- colors: 40, 40, 40, 40
			        1474 => x"00000000",		-- colors: 40, 40, 40, 40
			        1475 => x"00000000",		-- colors: 40, 40, 40, 40
			        1476 => x"00000000",		-- colors: 40, 40, 40, 40
			        1477 => x"00000000",		-- colors: 40, 40, 40, 40
			        1478 => x"00000000",		-- colors: 40, 40, 40, 40
			        1479 => x"00000000",		-- colors: 40, 40, 40, 40
			        1480 => x"00000000",		-- colors: 40, 40, 40, 40
			        1481 => x"00000000",		-- colors: 40, 40, 40, 40
			        1482 => x"00000000",		-- colors: 40, 40, 40, 40
			        1483 => x"00000000",		-- colors: 40, 40, 40, 40
			        1484 => x"00000000",		-- colors: 40, 40, 40, 40
			        1485 => x"00000000",		-- colors: 40, 40, 40, 40
			        1486 => x"00000000",		-- colors: 40, 40, 40, 40
			        1487 => x"00000000",		-- colors: 40, 40, 40, 40
			        1488 => x"00000000",		-- colors: 40, 40, 40, 40
			        1489 => x"00000000",		-- colors: 40, 40, 40, 40
			        1490 => x"00000000",		-- colors: 40, 40, 40, 40
			        1491 => x"00000000",		-- colors: 40, 40, 40, 40
			        1492 => x"00000000",		-- colors: 40, 40, 40, 40
			        1493 => x"00000000",		-- colors: 40, 40, 40, 40
			        1494 => x"00000000",		-- colors: 40, 40, 40, 40
			        1495 => x"00000000",		-- colors: 40, 40, 40, 40
			        1496 => x"00000000",		-- colors: 40, 40, 40, 40
			        1497 => x"00000000",		-- colors: 40, 40, 40, 40
			        1498 => x"00000000",		-- colors: 40, 40, 40, 40
			        1499 => x"00000000",		-- colors: 40, 40, 40, 40
			        1500 => x"00000000",		-- colors: 40, 40, 40, 40
			        1501 => x"00000000",		-- colors: 40, 40, 40, 40
			        1502 => x"00000000",		-- colors: 40, 40, 40, 40
			        1503 => x"00000000",		-- colors: 40, 40, 40, 40
			        1504 => x"00000000",		-- colors: 40, 40, 40, 40
			        1505 => x"00000000",		-- colors: 40, 40, 40, 40
			        1506 => x"00000000",		-- colors: 40, 40, 40, 40
			        1507 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1508 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1509 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1510 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1511 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1512 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1513 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1514 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1515 => x"00000000",		-- colors: 40, 40, 40, 40
			        1516 => x"00000000",		-- colors: 40, 40, 40, 40
			        1517 => x"00000000",		-- colors: 40, 40, 40, 40
			        1518 => x"00000000",		-- colors: 40, 40, 40, 40
			        1519 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1520 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1521 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1522 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1523 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1524 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1525 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1526 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1527 => x"00000000",		-- colors: 40, 40, 40, 40
			        1528 => x"00000000",		-- colors: 40, 40, 40, 40
			        1529 => x"00000000",		-- colors: 40, 40, 40, 40
			        1530 => x"00000000",		-- colors: 40, 40, 40, 40
			        1531 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1532 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1533 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1534 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60

			                --  sprite 20
			        1535 => x"00000000",		-- colors: 40, 40, 40, 40
			        1536 => x"00000000",		-- colors: 40, 40, 40, 40
			        1537 => x"00000000",		-- colors: 40, 40, 40, 40
			        1538 => x"00000000",		-- colors: 40, 40, 40, 40
			        1539 => x"00000000",		-- colors: 40, 40, 40, 40
			        1540 => x"00000000",		-- colors: 40, 40, 40, 40
			        1541 => x"00000000",		-- colors: 40, 40, 40, 40
			        1542 => x"00000000",		-- colors: 40, 40, 40, 40
			        1543 => x"00000000",		-- colors: 40, 40, 40, 40
			        1544 => x"00000000",		-- colors: 40, 40, 40, 40
			        1545 => x"00000000",		-- colors: 40, 40, 40, 40
			        1546 => x"00000000",		-- colors: 40, 40, 40, 40
			        1547 => x"00000000",		-- colors: 40, 40, 40, 40
			        1548 => x"00000000",		-- colors: 40, 40, 40, 40
			        1549 => x"00000000",		-- colors: 40, 40, 40, 40
			        1550 => x"00000000",		-- colors: 40, 40, 40, 40
			        1551 => x"00000000",		-- colors: 40, 40, 40, 40
			        1552 => x"00000000",		-- colors: 40, 40, 40, 40
			        1553 => x"00000000",		-- colors: 40, 40, 40, 40
			        1554 => x"00000000",		-- colors: 40, 40, 40, 40
			        1555 => x"00000000",		-- colors: 40, 40, 40, 40
			        1556 => x"00000000",		-- colors: 40, 40, 40, 40
			        1557 => x"00000000",		-- colors: 40, 40, 40, 40
			        1558 => x"00000000",		-- colors: 40, 40, 40, 40
			        1559 => x"00000000",		-- colors: 40, 40, 40, 40
			        1560 => x"00000000",		-- colors: 40, 40, 40, 40
			        1561 => x"00000000",		-- colors: 40, 40, 40, 40
			        1562 => x"00000000",		-- colors: 40, 40, 40, 40
			        1563 => x"00000000",		-- colors: 40, 40, 40, 40
			        1564 => x"00000000",		-- colors: 40, 40, 40, 40
			        1565 => x"00000000",		-- colors: 40, 40, 40, 40
			        1566 => x"00000000",		-- colors: 40, 40, 40, 40
			        1567 => x"00000000",		-- colors: 40, 40, 40, 40
			        1568 => x"00000000",		-- colors: 40, 40, 40, 40
			        1569 => x"00000000",		-- colors: 40, 40, 40, 40
			        1570 => x"00000000",		-- colors: 40, 40, 40, 40
			        1571 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1572 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1573 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1574 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1575 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1576 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1577 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1578 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1579 => x"00000000",		-- colors: 40, 40, 40, 40
			        1580 => x"00000000",		-- colors: 40, 40, 40, 40
			        1581 => x"00000000",		-- colors: 40, 40, 40, 40
			        1582 => x"00000000",		-- colors: 40, 40, 40, 40
			        1583 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1584 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1585 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1586 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1587 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1588 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1589 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1590 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1591 => x"00000000",		-- colors: 40, 40, 40, 40
			        1592 => x"00000000",		-- colors: 40, 40, 40, 40
			        1593 => x"00000000",		-- colors: 40, 40, 40, 40
			        1594 => x"00000000",		-- colors: 40, 40, 40, 40
			        1595 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1596 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1597 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1598 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60

			                --  sprite 21
			        1599 => x"3A3A3A3A",		-- colors: 58, 58, 58, 58
			        1600 => x"3A3A3A3A",		-- colors: 58, 58, 58, 58
			        1601 => x"3A3A3A3A",		-- colors: 58, 58, 58, 58
			        1602 => x"3A3A3A3A",		-- colors: 58, 58, 58, 58
			        1603 => x"3A3A3A3A",		-- colors: 58, 58, 58, 58
			        1604 => x"3A3A3A3A",		-- colors: 58, 58, 58, 58
			        1605 => x"3A3A3A3A",		-- colors: 58, 58, 58, 58
			        1606 => x"3A3A3A3A",		-- colors: 58, 58, 58, 58
			        1607 => x"3B3B3B3B",		-- colors: 59, 59, 59, 59
			        1608 => x"3B3B3B3B",		-- colors: 59, 59, 59, 59
			        1609 => x"3B3B3B3B",		-- colors: 59, 59, 59, 59
			        1610 => x"3B3B3B3B",		-- colors: 59, 59, 59, 59
			        1611 => x"39393939",		-- colors: 57, 57, 57, 57
			        1612 => x"39393939",		-- colors: 57, 57, 57, 57
			        1613 => x"39393939",		-- colors: 57, 57, 57, 57
			        1614 => x"39393939",		-- colors: 57, 57, 57, 57
			        1615 => x"39393939",		-- colors: 57, 57, 57, 57
			        1616 => x"39393939",		-- colors: 57, 57, 57, 57
			        1617 => x"39393939",		-- colors: 57, 57, 57, 57
			        1618 => x"39393939",		-- colors: 57, 57, 57, 57
			        1619 => x"39393939",		-- colors: 57, 57, 57, 57
			        1620 => x"39393939",		-- colors: 57, 57, 57, 57
			        1621 => x"39393939",		-- colors: 57, 57, 57, 57
			        1622 => x"39393939",		-- colors: 57, 57, 57, 57
			        1623 => x"39393939",		-- colors: 57, 57, 57, 57
			        1624 => x"39393939",		-- colors: 57, 57, 57, 57
			        1625 => x"39393939",		-- colors: 57, 57, 57, 57
			        1626 => x"39393939",		-- colors: 57, 57, 57, 57
			        1627 => x"39393939",		-- colors: 57, 57, 57, 57
			        1628 => x"39393939",		-- colors: 57, 57, 57, 57
			        1629 => x"39393939",		-- colors: 57, 57, 57, 57
			        1630 => x"39393939",		-- colors: 57, 57, 57, 57
			        1631 => x"39393939",		-- colors: 57, 57, 57, 57
			        1632 => x"39393939",		-- colors: 57, 57, 57, 57
			        1633 => x"39393939",		-- colors: 57, 57, 57, 57
			        1634 => x"39393939",		-- colors: 57, 57, 57, 57
			        1635 => x"39393939",		-- colors: 57, 57, 57, 57
			        1636 => x"39393939",		-- colors: 57, 57, 57, 57
			        1637 => x"39393939",		-- colors: 57, 57, 57, 57
			        1638 => x"39393939",		-- colors: 57, 57, 57, 57
			        1639 => x"39393939",		-- colors: 57, 57, 57, 57
			        1640 => x"39393939",		-- colors: 57, 57, 57, 57
			        1641 => x"39393939",		-- colors: 57, 57, 57, 57
			        1642 => x"39393939",		-- colors: 57, 57, 57, 57
			        1643 => x"39393939",		-- colors: 57, 57, 57, 57
			        1644 => x"39393939",		-- colors: 57, 57, 57, 57
			        1645 => x"39393939",		-- colors: 57, 57, 57, 57
			        1646 => x"39393939",		-- colors: 57, 57, 57, 57
			        1647 => x"39393939",		-- colors: 57, 57, 57, 57
			        1648 => x"39393939",		-- colors: 57, 57, 57, 57
			        1649 => x"39393939",		-- colors: 57, 57, 57, 57
			        1650 => x"39393939",		-- colors: 57, 57, 57, 57
			        1651 => x"39393939",		-- colors: 57, 57, 57, 57
			        1652 => x"39393939",		-- colors: 57, 57, 57, 57
			        1653 => x"39393939",		-- colors: 57, 57, 57, 57
			        1654 => x"39393939",		-- colors: 57, 57, 57, 57
			        1655 => x"39393939",		-- colors: 57, 57, 57, 57
			        1656 => x"39393939",		-- colors: 57, 57, 57, 57
			        1657 => x"39393939",		-- colors: 57, 57, 57, 57
			        1658 => x"39393939",		-- colors: 57, 57, 57, 57
			        1659 => x"3B3B3B3B",		-- colors: 59, 59, 59, 59
			        1660 => x"3B3B3B3B",		-- colors: 59, 59, 59, 59
			        1661 => x"3B3B3B3B",		-- colors: 59, 59, 59, 59
			        1662 => x"3B3B3B3B",		-- colors: 59, 59, 59, 59

			                --  sprite 22
			        1663 => x"00000000",		-- colors: 40, 40, 40, 40
			        1664 => x"00000000",		-- colors: 40, 40, 40, 40
			        1665 => x"00000000",		-- colors: 40, 40, 40, 40
			        1666 => x"00000000",		-- colors: 40, 40, 40, 40
			        1667 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1668 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1669 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1670 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1671 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1672 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1673 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1674 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1675 => x"00000000",		-- colors: 40, 40, 40, 40
			        1676 => x"00000000",		-- colors: 40, 40, 40, 40
			        1677 => x"00000000",		-- colors: 40, 40, 40, 40
			        1678 => x"00000000",		-- colors: 40, 40, 40, 40
			        1679 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1680 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1681 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1682 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1683 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1684 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1685 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1686 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1687 => x"00000000",		-- colors: 40, 40, 40, 40
			        1688 => x"00000000",		-- colors: 40, 40, 40, 40
			        1689 => x"00000000",		-- colors: 40, 40, 40, 40
			        1690 => x"00000000",		-- colors: 40, 40, 40, 40
			        1691 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1692 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1693 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1694 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1695 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1696 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1697 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1698 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1699 => x"00000000",		-- colors: 40, 40, 40, 40
			        1700 => x"00000000",		-- colors: 40, 40, 40, 40
			        1701 => x"00000000",		-- colors: 40, 40, 40, 40
			        1702 => x"00000000",		-- colors: 40, 40, 40, 40
			        1703 => x"00000000",		-- colors: 40, 40, 40, 40
			        1704 => x"00000000",		-- colors: 40, 40, 40, 40
			        1705 => x"00000000",		-- colors: 40, 40, 40, 40
			        1706 => x"00000000",		-- colors: 40, 40, 40, 40
			        1707 => x"00000000",		-- colors: 40, 40, 40, 40
			        1708 => x"00000000",		-- colors: 40, 40, 40, 40
			        1709 => x"00000000",		-- colors: 40, 40, 40, 40
			        1710 => x"00000000",		-- colors: 40, 40, 40, 40
			        1711 => x"00000000",		-- colors: 40, 40, 40, 40
			        1712 => x"00000000",		-- colors: 40, 40, 40, 40
			        1713 => x"00000000",		-- colors: 40, 40, 40, 40
			        1714 => x"00000000",		-- colors: 40, 40, 40, 40
			        1715 => x"00000000",		-- colors: 40, 40, 40, 40
			        1716 => x"00000000",		-- colors: 40, 40, 40, 40
			        1717 => x"00000000",		-- colors: 40, 40, 40, 40
			        1718 => x"00000000",		-- colors: 40, 40, 40, 40
			        1719 => x"00000000",		-- colors: 40, 40, 40, 40
			        1720 => x"00000000",		-- colors: 40, 40, 40, 40
			        1721 => x"00000000",		-- colors: 40, 40, 40, 40
			        1722 => x"00000000",		-- colors: 40, 40, 40, 40
			        1723 => x"00000000",		-- colors: 40, 40, 40, 40
			        1724 => x"00000000",		-- colors: 40, 40, 40, 40
			        1725 => x"00000000",		-- colors: 40, 40, 40, 40
			        1726 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 23
			        1727 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1728 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1729 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1730 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1731 => x"00000000",		-- colors: 40, 40, 40, 40
			        1732 => x"00000000",		-- colors: 40, 40, 40, 40
			        1733 => x"00000000",		-- colors: 40, 40, 40, 40
			        1734 => x"00000000",		-- colors: 40, 40, 40, 40
			        1735 => x"00000000",		-- colors: 40, 40, 40, 40
			        1736 => x"00000000",		-- colors: 40, 40, 40, 40
			        1737 => x"00000000",		-- colors: 40, 40, 40, 40
			        1738 => x"00000000",		-- colors: 40, 40, 40, 40
			        1739 => x"00000000",		-- colors: 40, 40, 40, 40
			        1740 => x"00000000",		-- colors: 40, 40, 40, 40
			        1741 => x"00000000",		-- colors: 40, 40, 40, 40
			        1742 => x"00000000",		-- colors: 40, 40, 40, 40
			        1743 => x"00000000",		-- colors: 40, 40, 40, 40
			        1744 => x"00000000",		-- colors: 40, 40, 40, 40
			        1745 => x"00000000",		-- colors: 40, 40, 40, 40
			        1746 => x"00000000",		-- colors: 40, 40, 40, 40
			        1747 => x"00000000",		-- colors: 40, 40, 40, 40
			        1748 => x"00000000",		-- colors: 40, 40, 40, 40
			        1749 => x"00000000",		-- colors: 40, 40, 40, 40
			        1750 => x"00000000",		-- colors: 40, 40, 40, 40
			        1751 => x"00000000",		-- colors: 40, 40, 40, 40
			        1752 => x"00000000",		-- colors: 40, 40, 40, 40
			        1753 => x"00000000",		-- colors: 40, 40, 40, 40
			        1754 => x"00000000",		-- colors: 40, 40, 40, 40
			        1755 => x"00000000",		-- colors: 40, 40, 40, 40
			        1756 => x"00000000",		-- colors: 40, 40, 40, 40
			        1757 => x"00000000",		-- colors: 40, 40, 40, 40
			        1758 => x"00000000",		-- colors: 40, 40, 40, 40
			        1759 => x"00000000",		-- colors: 40, 40, 40, 40
			        1760 => x"00000000",		-- colors: 40, 40, 40, 40
			        1761 => x"00000000",		-- colors: 40, 40, 40, 40
			        1762 => x"00000000",		-- colors: 40, 40, 40, 40
			        1763 => x"00000000",		-- colors: 40, 40, 40, 40
			        1764 => x"00000000",		-- colors: 40, 40, 40, 40
			        1765 => x"00000000",		-- colors: 40, 40, 40, 40
			        1766 => x"00000000",		-- colors: 40, 40, 40, 40
			        1767 => x"00000000",		-- colors: 40, 40, 40, 40
			        1768 => x"00000000",		-- colors: 40, 40, 40, 40
			        1769 => x"00000000",		-- colors: 40, 40, 40, 40
			        1770 => x"00000000",		-- colors: 40, 40, 40, 40
			        1771 => x"00000000",		-- colors: 40, 40, 40, 40
			        1772 => x"00000000",		-- colors: 40, 40, 40, 40
			        1773 => x"00000000",		-- colors: 40, 40, 40, 40
			        1774 => x"00000000",		-- colors: 40, 40, 40, 40
			        1775 => x"00000000",		-- colors: 40, 40, 40, 40
			        1776 => x"00000000",		-- colors: 40, 40, 40, 40
			        1777 => x"00000000",		-- colors: 40, 40, 40, 40
			        1778 => x"00000000",		-- colors: 40, 40, 40, 40
			        1779 => x"00000000",		-- colors: 40, 40, 40, 40
			        1780 => x"00000000",		-- colors: 40, 40, 40, 40
			        1781 => x"00000000",		-- colors: 40, 40, 40, 40
			        1782 => x"00000000",		-- colors: 40, 40, 40, 40
			        1783 => x"00000000",		-- colors: 40, 40, 40, 40
			        1784 => x"00000000",		-- colors: 40, 40, 40, 40
			        1785 => x"00000000",		-- colors: 40, 40, 40, 40
			        1786 => x"00000000",		-- colors: 40, 40, 40, 40
			        1787 => x"00000000",		-- colors: 40, 40, 40, 40
			        1788 => x"00000000",		-- colors: 40, 40, 40, 40
			        1789 => x"00000000",		-- colors: 40, 40, 40, 40
			        1790 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 24
			        1791 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1792 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1793 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1794 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1795 => x"00000000",		-- colors: 40, 40, 40, 40
			        1796 => x"00000000",		-- colors: 40, 40, 40, 40
			        1797 => x"00000000",		-- colors: 40, 40, 40, 40
			        1798 => x"00000000",		-- colors: 40, 40, 40, 40
			        1799 => x"00000000",		-- colors: 40, 40, 40, 40
			        1800 => x"00000000",		-- colors: 40, 40, 40, 40
			        1801 => x"00000000",		-- colors: 40, 40, 40, 40
			        1802 => x"00000000",		-- colors: 40, 40, 40, 40
			        1803 => x"00000000",		-- colors: 40, 40, 40, 40
			        1804 => x"00000000",		-- colors: 40, 40, 40, 40
			        1805 => x"00000000",		-- colors: 40, 40, 40, 40
			        1806 => x"00000000",		-- colors: 40, 40, 40, 40
			        1807 => x"00000000",		-- colors: 40, 40, 40, 40
			        1808 => x"00000000",		-- colors: 40, 40, 40, 40
			        1809 => x"00000000",		-- colors: 40, 40, 40, 40
			        1810 => x"00000000",		-- colors: 40, 40, 40, 40
			        1811 => x"00000000",		-- colors: 40, 40, 40, 40
			        1812 => x"00000000",		-- colors: 40, 40, 40, 40
			        1813 => x"00000000",		-- colors: 40, 40, 40, 40
			        1814 => x"00000000",		-- colors: 40, 40, 40, 40
			        1815 => x"00000000",		-- colors: 40, 40, 40, 40
			        1816 => x"00000000",		-- colors: 40, 40, 40, 40
			        1817 => x"00000000",		-- colors: 40, 40, 40, 40
			        1818 => x"00000000",		-- colors: 40, 40, 40, 40
			        1819 => x"00000000",		-- colors: 40, 40, 40, 40
			        1820 => x"00000000",		-- colors: 40, 40, 40, 40
			        1821 => x"00000000",		-- colors: 40, 40, 40, 40
			        1822 => x"00000000",		-- colors: 40, 40, 40, 40
			        1823 => x"00000000",		-- colors: 40, 40, 40, 40
			        1824 => x"00000000",		-- colors: 40, 40, 40, 40
			        1825 => x"00000000",		-- colors: 40, 40, 40, 40
			        1826 => x"00000000",		-- colors: 40, 40, 40, 40
			        1827 => x"00000000",		-- colors: 40, 40, 40, 40
			        1828 => x"00000000",		-- colors: 40, 40, 40, 40
			        1829 => x"00000000",		-- colors: 40, 40, 40, 40
			        1830 => x"00000000",		-- colors: 40, 40, 40, 40
			        1831 => x"00000000",		-- colors: 40, 40, 40, 40
			        1832 => x"00000000",		-- colors: 40, 40, 40, 40
			        1833 => x"00000000",		-- colors: 40, 40, 40, 40
			        1834 => x"00000000",		-- colors: 40, 40, 40, 40
			        1835 => x"00000000",		-- colors: 40, 40, 40, 40
			        1836 => x"00000000",		-- colors: 40, 40, 40, 40
			        1837 => x"00000000",		-- colors: 40, 40, 40, 40
			        1838 => x"00000000",		-- colors: 40, 40, 40, 40
			        1839 => x"00000000",		-- colors: 40, 40, 40, 40
			        1840 => x"00000000",		-- colors: 40, 40, 40, 40
			        1841 => x"00000000",		-- colors: 40, 40, 40, 40
			        1842 => x"00000000",		-- colors: 40, 40, 40, 40
			        1843 => x"00000000",		-- colors: 40, 40, 40, 40
			        1844 => x"00000000",		-- colors: 40, 40, 40, 40
			        1845 => x"00000000",		-- colors: 40, 40, 40, 40
			        1846 => x"00000000",		-- colors: 40, 40, 40, 40
			        1847 => x"00000000",		-- colors: 40, 40, 40, 40
			        1848 => x"00000000",		-- colors: 40, 40, 40, 40
			        1849 => x"00000000",		-- colors: 40, 40, 40, 40
			        1850 => x"00000000",		-- colors: 40, 40, 40, 40
			        1851 => x"00000000",		-- colors: 40, 40, 40, 40
			        1852 => x"00000000",		-- colors: 40, 40, 40, 40
			        1853 => x"00000000",		-- colors: 40, 40, 40, 40
			        1854 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 25
			        1855 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1856 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1857 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1858 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1859 => x"00000000",		-- colors: 40, 40, 40, 40
			        1860 => x"00000000",		-- colors: 40, 40, 40, 40
			        1861 => x"00000000",		-- colors: 40, 40, 40, 40
			        1862 => x"00000000",		-- colors: 40, 40, 40, 40
			        1863 => x"00000000",		-- colors: 40, 40, 40, 40
			        1864 => x"00000000",		-- colors: 40, 40, 40, 40
			        1865 => x"00000000",		-- colors: 40, 40, 40, 40
			        1866 => x"00000000",		-- colors: 40, 40, 40, 40
			        1867 => x"00000000",		-- colors: 40, 40, 40, 40
			        1868 => x"00000000",		-- colors: 40, 40, 40, 40
			        1869 => x"00000000",		-- colors: 40, 40, 40, 40
			        1870 => x"00000000",		-- colors: 40, 40, 40, 40
			        1871 => x"00000000",		-- colors: 40, 40, 40, 40
			        1872 => x"00000000",		-- colors: 40, 40, 40, 40
			        1873 => x"00000000",		-- colors: 40, 40, 40, 40
			        1874 => x"00000000",		-- colors: 40, 40, 40, 40
			        1875 => x"00000000",		-- colors: 40, 40, 40, 40
			        1876 => x"00000000",		-- colors: 40, 40, 40, 40
			        1877 => x"00000000",		-- colors: 40, 40, 40, 40
			        1878 => x"00000000",		-- colors: 40, 40, 40, 40
			        1879 => x"00000000",		-- colors: 40, 40, 40, 40
			        1880 => x"00000000",		-- colors: 40, 40, 40, 40
			        1881 => x"00000000",		-- colors: 40, 40, 40, 40
			        1882 => x"00000000",		-- colors: 40, 40, 40, 40
			        1883 => x"00000000",		-- colors: 40, 40, 40, 40
			        1884 => x"00000000",		-- colors: 40, 40, 40, 40
			        1885 => x"00000000",		-- colors: 40, 40, 40, 40
			        1886 => x"00000000",		-- colors: 40, 40, 40, 40
			        1887 => x"00000000",		-- colors: 40, 40, 40, 40
			        1888 => x"00000000",		-- colors: 40, 40, 40, 40
			        1889 => x"00000000",		-- colors: 40, 40, 40, 40
			        1890 => x"00000000",		-- colors: 40, 40, 40, 40
			        1891 => x"00000000",		-- colors: 40, 40, 40, 40
			        1892 => x"00000000",		-- colors: 40, 40, 40, 40
			        1893 => x"00000000",		-- colors: 40, 40, 40, 40
			        1894 => x"00000000",		-- colors: 40, 40, 40, 40
			        1895 => x"00000000",		-- colors: 40, 40, 40, 40
			        1896 => x"00000000",		-- colors: 40, 40, 40, 40
			        1897 => x"00000000",		-- colors: 40, 40, 40, 40
			        1898 => x"00000000",		-- colors: 40, 40, 40, 40
			        1899 => x"00000000",		-- colors: 40, 40, 40, 40
			        1900 => x"00000000",		-- colors: 40, 40, 40, 40
			        1901 => x"00000000",		-- colors: 40, 40, 40, 40
			        1902 => x"00000000",		-- colors: 40, 40, 40, 40
			        1903 => x"00000000",		-- colors: 40, 40, 40, 40
			        1904 => x"00000000",		-- colors: 40, 40, 40, 40
			        1905 => x"00000000",		-- colors: 40, 40, 40, 40
			        1906 => x"00000000",		-- colors: 40, 40, 40, 40
			        1907 => x"00000000",		-- colors: 40, 40, 40, 40
			        1908 => x"00000000",		-- colors: 40, 40, 40, 40
			        1909 => x"00000000",		-- colors: 40, 40, 40, 40
			        1910 => x"00000000",		-- colors: 40, 40, 40, 40
			        1911 => x"00000000",		-- colors: 40, 40, 40, 40
			        1912 => x"00000000",		-- colors: 40, 40, 40, 40
			        1913 => x"00000000",		-- colors: 40, 40, 40, 40
			        1914 => x"00000000",		-- colors: 40, 40, 40, 40
			        1915 => x"00000000",		-- colors: 40, 40, 40, 40
			        1916 => x"00000000",		-- colors: 40, 40, 40, 40
			        1917 => x"00000000",		-- colors: 40, 40, 40, 40
			        1918 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 26
			        1919 => x"3A3A3A3A",		-- colors: 58, 58, 58, 58
			        1920 => x"3A3A3A3A",		-- colors: 58, 58, 58, 58
			        1921 => x"3A3A3A3A",		-- colors: 58, 58, 58, 58
			        1922 => x"3A3A3A3A",		-- colors: 58, 58, 58, 58
			        1923 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1924 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1925 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1926 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1927 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1928 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1929 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1930 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1931 => x"00000000",		-- colors: 40, 40, 40, 40
			        1932 => x"00000000",		-- colors: 40, 40, 40, 40
			        1933 => x"00000000",		-- colors: 40, 40, 40, 40
			        1934 => x"00000000",		-- colors: 40, 40, 40, 40
			        1935 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1936 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1937 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1938 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1939 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1940 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1941 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1942 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1943 => x"00000000",		-- colors: 40, 40, 40, 40
			        1944 => x"00000000",		-- colors: 40, 40, 40, 40
			        1945 => x"00000000",		-- colors: 40, 40, 40, 40
			        1946 => x"00000000",		-- colors: 40, 40, 40, 40
			        1947 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1948 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1949 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1950 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1951 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1952 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1953 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1954 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1955 => x"00000000",		-- colors: 40, 40, 40, 40
			        1956 => x"00000000",		-- colors: 40, 40, 40, 40
			        1957 => x"00000000",		-- colors: 40, 40, 40, 40
			        1958 => x"00000000",		-- colors: 40, 40, 40, 40
			        1959 => x"00000000",		-- colors: 40, 40, 40, 40
			        1960 => x"00000000",		-- colors: 40, 40, 40, 40
			        1961 => x"00000000",		-- colors: 40, 40, 40, 40
			        1962 => x"00000000",		-- colors: 40, 40, 40, 40
			        1963 => x"00000000",		-- colors: 40, 40, 40, 40
			        1964 => x"00000000",		-- colors: 40, 40, 40, 40
			        1965 => x"00000000",		-- colors: 40, 40, 40, 40
			        1966 => x"00000000",		-- colors: 40, 40, 40, 40
			        1967 => x"00000000",		-- colors: 40, 40, 40, 40
			        1968 => x"00000000",		-- colors: 40, 40, 40, 40
			        1969 => x"00000000",		-- colors: 40, 40, 40, 40
			        1970 => x"00000000",		-- colors: 40, 40, 40, 40
			        1971 => x"00000000",		-- colors: 40, 40, 40, 40
			        1972 => x"00000000",		-- colors: 40, 40, 40, 40
			        1973 => x"00000000",		-- colors: 40, 40, 40, 40
			        1974 => x"00000000",		-- colors: 40, 40, 40, 40
			        1975 => x"00000000",		-- colors: 40, 40, 40, 40
			        1976 => x"00000000",		-- colors: 40, 40, 40, 40
			        1977 => x"00000000",		-- colors: 40, 40, 40, 40
			        1978 => x"00000000",		-- colors: 40, 40, 40, 40
			        1979 => x"00000000",		-- colors: 40, 40, 40, 40
			        1980 => x"00000000",		-- colors: 40, 40, 40, 40
			        1981 => x"00000000",		-- colors: 40, 40, 40, 40
			        1982 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 27
			        1983 => x"00000000",		-- colors: 40, 40, 40, 40
			        1984 => x"00000000",		-- colors: 40, 40, 40, 40
			        1985 => x"00000000",		-- colors: 40, 40, 40, 40
			        1986 => x"00000000",		-- colors: 40, 40, 40, 40
			        1987 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1988 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1989 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1990 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1991 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1992 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1993 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1994 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        1995 => x"00000000",		-- colors: 40, 40, 40, 40
			        1996 => x"00000000",		-- colors: 40, 40, 40, 40
			        1997 => x"00000000",		-- colors: 40, 40, 40, 40
			        1998 => x"00000000",		-- colors: 40, 40, 40, 40
			        1999 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2000 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2001 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2002 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2003 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2004 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2005 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2006 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2007 => x"00000000",		-- colors: 40, 40, 40, 40
			        2008 => x"00000000",		-- colors: 40, 40, 40, 40
			        2009 => x"00000000",		-- colors: 40, 40, 40, 40
			        2010 => x"00000000",		-- colors: 40, 40, 40, 40
			        2011 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2012 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2013 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2014 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2015 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2016 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2017 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2018 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2019 => x"00000000",		-- colors: 40, 40, 40, 40
			        2020 => x"00000000",		-- colors: 40, 40, 40, 40
			        2021 => x"00000000",		-- colors: 40, 40, 40, 40
			        2022 => x"00000000",		-- colors: 40, 40, 40, 40
			        2023 => x"00000000",		-- colors: 40, 40, 40, 40
			        2024 => x"00000000",		-- colors: 40, 40, 40, 40
			        2025 => x"00000000",		-- colors: 40, 40, 40, 40
			        2026 => x"00000000",		-- colors: 40, 40, 40, 40
			        2027 => x"00000000",		-- colors: 40, 40, 40, 40
			        2028 => x"00000000",		-- colors: 40, 40, 40, 40
			        2029 => x"00000000",		-- colors: 40, 40, 40, 40
			        2030 => x"00000000",		-- colors: 40, 40, 40, 40
			        2031 => x"00000000",		-- colors: 40, 40, 40, 40
			        2032 => x"00000000",		-- colors: 40, 40, 40, 40
			        2033 => x"00000000",		-- colors: 40, 40, 40, 40
			        2034 => x"00000000",		-- colors: 40, 40, 40, 40
			        2035 => x"00000000",		-- colors: 40, 40, 40, 40
			        2036 => x"00000000",		-- colors: 40, 40, 40, 40
			        2037 => x"00000000",		-- colors: 40, 40, 40, 40
			        2038 => x"00000000",		-- colors: 40, 40, 40, 40
			        2039 => x"00000000",		-- colors: 40, 40, 40, 40
			        2040 => x"00000000",		-- colors: 40, 40, 40, 40
			        2041 => x"00000000",		-- colors: 40, 40, 40, 40
			        2042 => x"00000000",		-- colors: 40, 40, 40, 40
			        2043 => x"00000000",		-- colors: 40, 40, 40, 40
			        2044 => x"00000000",		-- colors: 40, 40, 40, 40
			        2045 => x"00000000",		-- colors: 40, 40, 40, 40
			        2046 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 28
			        2047 => x"00000000",		-- colors: 40, 40, 40, 40
			        2048 => x"00000000",		-- colors: 40, 40, 40, 40
			        2049 => x"00000000",		-- colors: 40, 40, 40, 40
			        2050 => x"00000000",		-- colors: 40, 40, 40, 40
			        2051 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2052 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2053 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2054 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2055 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2056 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2057 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2058 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2059 => x"00000000",		-- colors: 40, 40, 40, 40
			        2060 => x"00000000",		-- colors: 40, 40, 40, 40
			        2061 => x"00000000",		-- colors: 40, 40, 40, 40
			        2062 => x"00000000",		-- colors: 40, 40, 40, 40
			        2063 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2064 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2065 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2066 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2067 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2068 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2069 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2070 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2071 => x"00000000",		-- colors: 40, 40, 40, 40
			        2072 => x"00000000",		-- colors: 40, 40, 40, 40
			        2073 => x"00000000",		-- colors: 40, 40, 40, 40
			        2074 => x"00000000",		-- colors: 40, 40, 40, 40
			        2075 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2076 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2077 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2078 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2079 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2080 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2081 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2082 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2083 => x"00000000",		-- colors: 40, 40, 40, 40
			        2084 => x"00000000",		-- colors: 40, 40, 40, 40
			        2085 => x"00000000",		-- colors: 40, 40, 40, 40
			        2086 => x"00000000",		-- colors: 40, 40, 40, 40
			        2087 => x"00000000",		-- colors: 40, 40, 40, 40
			        2088 => x"00000000",		-- colors: 40, 40, 40, 40
			        2089 => x"00000000",		-- colors: 40, 40, 40, 40
			        2090 => x"00000000",		-- colors: 40, 40, 40, 40
			        2091 => x"00000000",		-- colors: 40, 40, 40, 40
			        2092 => x"00000000",		-- colors: 40, 40, 40, 40
			        2093 => x"00000000",		-- colors: 40, 40, 40, 40
			        2094 => x"00000000",		-- colors: 40, 40, 40, 40
			        2095 => x"00000000",		-- colors: 40, 40, 40, 40
			        2096 => x"00000000",		-- colors: 40, 40, 40, 40
			        2097 => x"00000000",		-- colors: 40, 40, 40, 40
			        2098 => x"00000000",		-- colors: 40, 40, 40, 40
			        2099 => x"00000000",		-- colors: 40, 40, 40, 40
			        2100 => x"00000000",		-- colors: 40, 40, 40, 40
			        2101 => x"00000000",		-- colors: 40, 40, 40, 40
			        2102 => x"00000000",		-- colors: 40, 40, 40, 40
			        2103 => x"00000000",		-- colors: 40, 40, 40, 40
			        2104 => x"00000000",		-- colors: 40, 40, 40, 40
			        2105 => x"00000000",		-- colors: 40, 40, 40, 40
			        2106 => x"00000000",		-- colors: 40, 40, 40, 40
			        2107 => x"00000000",		-- colors: 40, 40, 40, 40
			        2108 => x"00000000",		-- colors: 40, 40, 40, 40
			        2109 => x"00000000",		-- colors: 40, 40, 40, 40
			        2110 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 29
			        2111 => x"00000000",		-- colors: 40, 40, 40, 40
			        2112 => x"00000000",		-- colors: 40, 40, 40, 40
			        2113 => x"00000000",		-- colors: 40, 40, 40, 40
			        2114 => x"00000000",		-- colors: 40, 40, 40, 40
			        2115 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2116 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2117 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2118 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2119 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2120 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2121 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2122 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2123 => x"00000000",		-- colors: 40, 40, 40, 40
			        2124 => x"00000000",		-- colors: 40, 40, 40, 40
			        2125 => x"00000000",		-- colors: 40, 40, 40, 40
			        2126 => x"00000000",		-- colors: 40, 40, 40, 40
			        2127 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2128 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2129 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2130 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2131 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2132 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2133 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2134 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2135 => x"00000000",		-- colors: 40, 40, 40, 40
			        2136 => x"00000000",		-- colors: 40, 40, 40, 40
			        2137 => x"00000000",		-- colors: 40, 40, 40, 40
			        2138 => x"00000000",		-- colors: 40, 40, 40, 40
			        2139 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2140 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2141 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2142 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2143 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2144 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2145 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2146 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2147 => x"00000000",		-- colors: 40, 40, 40, 40
			        2148 => x"00000000",		-- colors: 40, 40, 40, 40
			        2149 => x"00000000",		-- colors: 40, 40, 40, 40
			        2150 => x"00000000",		-- colors: 40, 40, 40, 40
			        2151 => x"00000000",		-- colors: 40, 40, 40, 40
			        2152 => x"00000000",		-- colors: 40, 40, 40, 40
			        2153 => x"00000000",		-- colors: 40, 40, 40, 40
			        2154 => x"00000000",		-- colors: 40, 40, 40, 40
			        2155 => x"00000000",		-- colors: 40, 40, 40, 40
			        2156 => x"00000000",		-- colors: 40, 40, 40, 40
			        2157 => x"00000000",		-- colors: 40, 40, 40, 40
			        2158 => x"00000000",		-- colors: 40, 40, 40, 40
			        2159 => x"00000000",		-- colors: 40, 40, 40, 40
			        2160 => x"00000000",		-- colors: 40, 40, 40, 40
			        2161 => x"00000000",		-- colors: 40, 40, 40, 40
			        2162 => x"00000000",		-- colors: 40, 40, 40, 40
			        2163 => x"00000000",		-- colors: 40, 40, 40, 40
			        2164 => x"00000000",		-- colors: 40, 40, 40, 40
			        2165 => x"00000000",		-- colors: 40, 40, 40, 40
			        2166 => x"00000000",		-- colors: 40, 40, 40, 40
			        2167 => x"00000000",		-- colors: 40, 40, 40, 40
			        2168 => x"00000000",		-- colors: 40, 40, 40, 40
			        2169 => x"00000000",		-- colors: 40, 40, 40, 40
			        2170 => x"00000000",		-- colors: 40, 40, 40, 40
			        2171 => x"00000000",		-- colors: 40, 40, 40, 40
			        2172 => x"00000000",		-- colors: 40, 40, 40, 40
			        2173 => x"00000000",		-- colors: 40, 40, 40, 40
			        2174 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 30
			        2175 => x"00000000",		-- colors: 40, 40, 40, 40
			        2176 => x"00000000",		-- colors: 40, 40, 40, 40
			        2177 => x"00000000",		-- colors: 40, 40, 40, 40
			        2178 => x"00000000",		-- colors: 40, 40, 40, 40
			        2179 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2180 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2181 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2182 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2183 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2184 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2185 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2186 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2187 => x"00000000",		-- colors: 40, 40, 40, 40
			        2188 => x"00000000",		-- colors: 40, 40, 40, 40
			        2189 => x"00000000",		-- colors: 40, 40, 40, 40
			        2190 => x"00000000",		-- colors: 40, 40, 40, 40
			        2191 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2192 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2193 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2194 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2195 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2196 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2197 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2198 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2199 => x"00000000",		-- colors: 40, 40, 40, 40
			        2200 => x"00000000",		-- colors: 40, 40, 40, 40
			        2201 => x"00000000",		-- colors: 40, 40, 40, 40
			        2202 => x"00000000",		-- colors: 40, 40, 40, 40
			        2203 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2204 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2205 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2206 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2207 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2208 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2209 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2210 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2211 => x"00000000",		-- colors: 40, 40, 40, 40
			        2212 => x"00000000",		-- colors: 40, 40, 40, 40
			        2213 => x"00000000",		-- colors: 40, 40, 40, 40
			        2214 => x"00000000",		-- colors: 40, 40, 40, 40
			        2215 => x"00000000",		-- colors: 40, 40, 40, 40
			        2216 => x"00000000",		-- colors: 40, 40, 40, 40
			        2217 => x"00000000",		-- colors: 40, 40, 40, 40
			        2218 => x"00000000",		-- colors: 40, 40, 40, 40
			        2219 => x"00000000",		-- colors: 40, 40, 40, 40
			        2220 => x"00000000",		-- colors: 40, 40, 40, 40
			        2221 => x"00000000",		-- colors: 40, 40, 40, 40
			        2222 => x"00000000",		-- colors: 40, 40, 40, 40
			        2223 => x"00000000",		-- colors: 40, 40, 40, 40
			        2224 => x"00000000",		-- colors: 40, 40, 40, 40
			        2225 => x"00000000",		-- colors: 40, 40, 40, 40
			        2226 => x"00000000",		-- colors: 40, 40, 40, 40
			        2227 => x"00000000",		-- colors: 40, 40, 40, 40
			        2228 => x"00000000",		-- colors: 40, 40, 40, 40
			        2229 => x"00000000",		-- colors: 40, 40, 40, 40
			        2230 => x"00000000",		-- colors: 40, 40, 40, 40
			        2231 => x"00000000",		-- colors: 40, 40, 40, 40
			        2232 => x"00000000",		-- colors: 40, 40, 40, 40
			        2233 => x"00000000",		-- colors: 40, 40, 40, 40
			        2234 => x"00000000",		-- colors: 40, 40, 40, 40
			        2235 => x"00000000",		-- colors: 40, 40, 40, 40
			        2236 => x"00000000",		-- colors: 40, 40, 40, 40
			        2237 => x"00000000",		-- colors: 40, 40, 40, 40
			        2238 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 31
			        2239 => x"00000000",		-- colors: 40, 40, 40, 40
			        2240 => x"00000000",		-- colors: 40, 40, 40, 40
			        2241 => x"00000000",		-- colors: 40, 40, 40, 40
			        2242 => x"00000000",		-- colors: 40, 40, 40, 40
			        2243 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2244 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2245 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2246 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2247 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2248 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2249 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2250 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2251 => x"00000000",		-- colors: 40, 40, 40, 40
			        2252 => x"00000000",		-- colors: 40, 40, 40, 40
			        2253 => x"00000000",		-- colors: 40, 40, 40, 40
			        2254 => x"00000000",		-- colors: 40, 40, 40, 40
			        2255 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2256 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2257 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2258 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2259 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2260 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2261 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2262 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2263 => x"00000000",		-- colors: 40, 40, 40, 40
			        2264 => x"00000000",		-- colors: 40, 40, 40, 40
			        2265 => x"00000000",		-- colors: 40, 40, 40, 40
			        2266 => x"00000000",		-- colors: 40, 40, 40, 40
			        2267 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2268 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2269 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2270 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2271 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2272 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2273 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2274 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2275 => x"00000000",		-- colors: 40, 40, 40, 40
			        2276 => x"00000000",		-- colors: 40, 40, 40, 40
			        2277 => x"00000000",		-- colors: 40, 40, 40, 40
			        2278 => x"00000000",		-- colors: 40, 40, 40, 40
			        2279 => x"32323232",		-- colors: 50, 50, 50, 50
			        2280 => x"32323232",		-- colors: 50, 50, 50, 50
			        2281 => x"32323232",		-- colors: 50, 50, 50, 50
			        2282 => x"32323232",		-- colors: 50, 50, 50, 50
			        2283 => x"00000000",		-- colors: 40, 40, 40, 40
			        2284 => x"00000000",		-- colors: 40, 40, 40, 40
			        2285 => x"00000000",		-- colors: 40, 40, 40, 40
			        2286 => x"00000000",		-- colors: 40, 40, 40, 40
			        2287 => x"00000000",		-- colors: 40, 40, 40, 40
			        2288 => x"00000000",		-- colors: 40, 40, 40, 40
			        2289 => x"00000000",		-- colors: 40, 40, 40, 40
			        2290 => x"00000000",		-- colors: 40, 40, 40, 40
			        2291 => x"00000000",		-- colors: 40, 40, 40, 40
			        2292 => x"00000000",		-- colors: 40, 40, 40, 40
			        2293 => x"00000000",		-- colors: 40, 40, 40, 40
			        2294 => x"00000000",		-- colors: 40, 40, 40, 40
			        2295 => x"32323232",		-- colors: 50, 50, 50, 50
			        2296 => x"32323232",		-- colors: 50, 50, 50, 50
			        2297 => x"32323232",		-- colors: 50, 50, 50, 50
			        2298 => x"32323232",		-- colors: 50, 50, 50, 50
			        2299 => x"00000000",		-- colors: 40, 40, 40, 40
			        2300 => x"00000000",		-- colors: 40, 40, 40, 40
			        2301 => x"00000000",		-- colors: 40, 40, 40, 40
			        2302 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 32
			        2303 => x"00000000",		-- colors: 40, 40, 40, 40
			        2304 => x"00000000",		-- colors: 40, 40, 40, 40
			        2305 => x"00000000",		-- colors: 40, 40, 40, 40
			        2306 => x"00000000",		-- colors: 40, 40, 40, 40
			        2307 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2308 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2309 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2310 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2311 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2312 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2313 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2314 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2315 => x"00000000",		-- colors: 40, 40, 40, 40
			        2316 => x"00000000",		-- colors: 40, 40, 40, 40
			        2317 => x"00000000",		-- colors: 40, 40, 40, 40
			        2318 => x"00000000",		-- colors: 40, 40, 40, 40
			        2319 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2320 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2321 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2322 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2323 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2324 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2325 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2326 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2327 => x"00000000",		-- colors: 40, 40, 40, 40
			        2328 => x"00000000",		-- colors: 40, 40, 40, 40
			        2329 => x"00000000",		-- colors: 40, 40, 40, 40
			        2330 => x"00000000",		-- colors: 40, 40, 40, 40
			        2331 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2332 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2333 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2334 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2335 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2336 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2337 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2338 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2339 => x"00000000",		-- colors: 40, 40, 40, 40
			        2340 => x"00000000",		-- colors: 40, 40, 40, 40
			        2341 => x"00000000",		-- colors: 40, 40, 40, 40
			        2342 => x"00000000",		-- colors: 40, 40, 40, 40
			        2343 => x"00000000",		-- colors: 40, 40, 40, 40
			        2344 => x"00000000",		-- colors: 40, 40, 40, 40
			        2345 => x"00000000",		-- colors: 40, 40, 40, 40
			        2346 => x"00000000",		-- colors: 40, 40, 40, 40
			        2347 => x"00000000",		-- colors: 40, 40, 40, 40
			        2348 => x"00000000",		-- colors: 40, 40, 40, 40
			        2349 => x"00000000",		-- colors: 40, 40, 40, 40
			        2350 => x"00000000",		-- colors: 40, 40, 40, 40
			        2351 => x"00000000",		-- colors: 40, 40, 40, 40
			        2352 => x"00000000",		-- colors: 40, 40, 40, 40
			        2353 => x"00000000",		-- colors: 40, 40, 40, 40
			        2354 => x"00000000",		-- colors: 40, 40, 40, 40
			        2355 => x"00000000",		-- colors: 40, 40, 40, 40
			        2356 => x"00000000",		-- colors: 40, 40, 40, 40
			        2357 => x"00000000",		-- colors: 40, 40, 40, 40
			        2358 => x"00000000",		-- colors: 40, 40, 40, 40
			        2359 => x"00000000",		-- colors: 40, 40, 40, 40
			        2360 => x"00000000",		-- colors: 40, 40, 40, 40
			        2361 => x"00000000",		-- colors: 40, 40, 40, 40
			        2362 => x"00000000",		-- colors: 40, 40, 40, 40
			        2363 => x"00000000",		-- colors: 40, 40, 40, 40
			        2364 => x"00000000",		-- colors: 40, 40, 40, 40
			        2365 => x"00000000",		-- colors: 40, 40, 40, 40
			        2366 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 33
			        2367 => x"00000000",		-- colors: 40, 40, 40, 40
			        2368 => x"00000000",		-- colors: 40, 40, 40, 40
			        2369 => x"00000000",		-- colors: 40, 40, 40, 40
			        2370 => x"00000000",		-- colors: 40, 40, 40, 40
			        2371 => x"00000000",		-- colors: 40, 40, 40, 40
			        2372 => x"00000000",		-- colors: 40, 40, 40, 40
			        2373 => x"00000000",		-- colors: 40, 40, 40, 40
			        2374 => x"00000000",		-- colors: 40, 40, 40, 40
			        2375 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2376 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2377 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2378 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2379 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2380 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2381 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2382 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2383 => x"00000000",		-- colors: 40, 40, 40, 40
			        2384 => x"00000000",		-- colors: 40, 40, 40, 40
			        2385 => x"00000000",		-- colors: 40, 40, 40, 40
			        2386 => x"00000000",		-- colors: 40, 40, 40, 40
			        2387 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2388 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2389 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2390 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2391 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2392 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2393 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2394 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2395 => x"00000000",		-- colors: 40, 40, 40, 40
			        2396 => x"00000000",		-- colors: 40, 40, 40, 40
			        2397 => x"00000000",		-- colors: 40, 40, 40, 40
			        2398 => x"00000000",		-- colors: 40, 40, 40, 40
			        2399 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2400 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2401 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2402 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2403 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2404 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2405 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2406 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2407 => x"00000000",		-- colors: 40, 40, 40, 40
			        2408 => x"00000000",		-- colors: 40, 40, 40, 40
			        2409 => x"00000000",		-- colors: 40, 40, 40, 40
			        2410 => x"00000000",		-- colors: 40, 40, 40, 40
			        2411 => x"00000000",		-- colors: 40, 40, 40, 40
			        2412 => x"00000000",		-- colors: 40, 40, 40, 40
			        2413 => x"00000000",		-- colors: 40, 40, 40, 40
			        2414 => x"00000000",		-- colors: 40, 40, 40, 40
			        2415 => x"00000000",		-- colors: 40, 40, 40, 40
			        2416 => x"00000000",		-- colors: 40, 40, 40, 40
			        2417 => x"00000000",		-- colors: 40, 40, 40, 40
			        2418 => x"00000000",		-- colors: 40, 40, 40, 40
			        2419 => x"00000000",		-- colors: 40, 40, 40, 40
			        2420 => x"00000000",		-- colors: 40, 40, 40, 40
			        2421 => x"00000000",		-- colors: 40, 40, 40, 40
			        2422 => x"00000000",		-- colors: 40, 40, 40, 40
			        2423 => x"00000000",		-- colors: 40, 40, 40, 40
			        2424 => x"00000000",		-- colors: 40, 40, 40, 40
			        2425 => x"00000000",		-- colors: 40, 40, 40, 40
			        2426 => x"00000000",		-- colors: 40, 40, 40, 40
			        2427 => x"00000000",		-- colors: 40, 40, 40, 40
			        2428 => x"00000000",		-- colors: 40, 40, 40, 40
			        2429 => x"00000000",		-- colors: 40, 40, 40, 40
			        2430 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 34
			        2431 => x"00000000",		-- colors: 40, 40, 40, 40
			        2432 => x"00000000",		-- colors: 40, 40, 40, 40
			        2433 => x"00000000",		-- colors: 40, 40, 40, 40
			        2434 => x"00000000",		-- colors: 40, 40, 40, 40
			        2435 => x"00000000",		-- colors: 40, 40, 40, 40
			        2436 => x"00000000",		-- colors: 40, 40, 40, 40
			        2437 => x"00000000",		-- colors: 40, 40, 40, 40
			        2438 => x"00000000",		-- colors: 40, 40, 40, 40
			        2439 => x"00000000",		-- colors: 40, 40, 40, 40
			        2440 => x"00000000",		-- colors: 40, 40, 40, 40
			        2441 => x"00000000",		-- colors: 40, 40, 40, 40
			        2442 => x"00000000",		-- colors: 40, 40, 40, 40
			        2443 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2444 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2445 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2446 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2447 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2448 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2449 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2450 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2451 => x"00000000",		-- colors: 40, 40, 40, 40
			        2452 => x"00000000",		-- colors: 40, 40, 40, 40
			        2453 => x"00000000",		-- colors: 40, 40, 40, 40
			        2454 => x"00000000",		-- colors: 40, 40, 40, 40
			        2455 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2456 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2457 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2458 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2459 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2460 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2461 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2462 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2463 => x"00000000",		-- colors: 40, 40, 40, 40
			        2464 => x"00000000",		-- colors: 40, 40, 40, 40
			        2465 => x"00000000",		-- colors: 40, 40, 40, 40
			        2466 => x"00000000",		-- colors: 40, 40, 40, 40
			        2467 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2468 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2469 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2470 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2471 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2472 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2473 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2474 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2475 => x"00000000",		-- colors: 40, 40, 40, 40
			        2476 => x"00000000",		-- colors: 40, 40, 40, 40
			        2477 => x"00000000",		-- colors: 40, 40, 40, 40
			        2478 => x"00000000",		-- colors: 40, 40, 40, 40
			        2479 => x"00000000",		-- colors: 40, 40, 40, 40
			        2480 => x"00000000",		-- colors: 40, 40, 40, 40
			        2481 => x"00000000",		-- colors: 40, 40, 40, 40
			        2482 => x"00000000",		-- colors: 40, 40, 40, 40
			        2483 => x"00000000",		-- colors: 40, 40, 40, 40
			        2484 => x"00000000",		-- colors: 40, 40, 40, 40
			        2485 => x"00000000",		-- colors: 40, 40, 40, 40
			        2486 => x"00000000",		-- colors: 40, 40, 40, 40
			        2487 => x"00000000",		-- colors: 40, 40, 40, 40
			        2488 => x"00000000",		-- colors: 40, 40, 40, 40
			        2489 => x"00000000",		-- colors: 40, 40, 40, 40
			        2490 => x"00000000",		-- colors: 40, 40, 40, 40
			        2491 => x"00000000",		-- colors: 40, 40, 40, 40
			        2492 => x"00000000",		-- colors: 40, 40, 40, 40
			        2493 => x"00000000",		-- colors: 40, 40, 40, 40
			        2494 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 35
			        2495 => x"00000000",		-- colors: 40, 40, 40, 40
			        2496 => x"00000000",		-- colors: 40, 40, 40, 40
			        2497 => x"00000000",		-- colors: 40, 40, 40, 40
			        2498 => x"00000000",		-- colors: 40, 40, 40, 40
			        2499 => x"00000000",		-- colors: 40, 40, 40, 40
			        2500 => x"00000000",		-- colors: 40, 40, 40, 40
			        2501 => x"00000000",		-- colors: 40, 40, 40, 40
			        2502 => x"00000000",		-- colors: 40, 40, 40, 40
			        2503 => x"00000000",		-- colors: 40, 40, 40, 40
			        2504 => x"00000000",		-- colors: 40, 40, 40, 40
			        2505 => x"00000000",		-- colors: 40, 40, 40, 40
			        2506 => x"00000000",		-- colors: 40, 40, 40, 40
			        2507 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2508 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2509 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2510 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2511 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2512 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2513 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2514 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2515 => x"00000000",		-- colors: 40, 40, 40, 40
			        2516 => x"00000000",		-- colors: 40, 40, 40, 40
			        2517 => x"00000000",		-- colors: 40, 40, 40, 40
			        2518 => x"00000000",		-- colors: 40, 40, 40, 40
			        2519 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2520 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2521 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2522 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2523 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2524 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2525 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2526 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2527 => x"00000000",		-- colors: 40, 40, 40, 40
			        2528 => x"00000000",		-- colors: 40, 40, 40, 40
			        2529 => x"00000000",		-- colors: 40, 40, 40, 40
			        2530 => x"00000000",		-- colors: 40, 40, 40, 40
			        2531 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2532 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2533 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2534 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2535 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2536 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2537 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2538 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2539 => x"00000000",		-- colors: 40, 40, 40, 40
			        2540 => x"00000000",		-- colors: 40, 40, 40, 40
			        2541 => x"00000000",		-- colors: 40, 40, 40, 40
			        2542 => x"00000000",		-- colors: 40, 40, 40, 40
			        2543 => x"00000000",		-- colors: 40, 40, 40, 40
			        2544 => x"00000000",		-- colors: 40, 40, 40, 40
			        2545 => x"00000000",		-- colors: 40, 40, 40, 40
			        2546 => x"00000000",		-- colors: 40, 40, 40, 40
			        2547 => x"00000000",		-- colors: 40, 40, 40, 40
			        2548 => x"00000000",		-- colors: 40, 40, 40, 40
			        2549 => x"00000000",		-- colors: 40, 40, 40, 40
			        2550 => x"00000000",		-- colors: 40, 40, 40, 40
			        2551 => x"00000000",		-- colors: 40, 40, 40, 40
			        2552 => x"00000000",		-- colors: 40, 40, 40, 40
			        2553 => x"00000000",		-- colors: 40, 40, 40, 40
			        2554 => x"00000000",		-- colors: 40, 40, 40, 40
			        2555 => x"00000000",		-- colors: 40, 40, 40, 40
			        2556 => x"00000000",		-- colors: 40, 40, 40, 40
			        2557 => x"00000000",		-- colors: 40, 40, 40, 40
			        2558 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 36
			        2559 => x"00000000",		-- colors: 40, 40, 40, 40
			        2560 => x"00000000",		-- colors: 40, 40, 40, 40
			        2561 => x"00000000",		-- colors: 40, 40, 40, 40
			        2562 => x"00000000",		-- colors: 40, 40, 40, 40
			        2563 => x"00000000",		-- colors: 40, 40, 40, 40
			        2564 => x"00000000",		-- colors: 40, 40, 40, 40
			        2565 => x"00000000",		-- colors: 40, 40, 40, 40
			        2566 => x"00000000",		-- colors: 40, 40, 40, 40
			        2567 => x"00000000",		-- colors: 40, 40, 40, 40
			        2568 => x"00000000",		-- colors: 40, 40, 40, 40
			        2569 => x"00000000",		-- colors: 40, 40, 40, 40
			        2570 => x"00000000",		-- colors: 40, 40, 40, 40
			        2571 => x"00000000",		-- colors: 40, 40, 40, 40
			        2572 => x"00000000",		-- colors: 40, 40, 40, 40
			        2573 => x"00000000",		-- colors: 40, 40, 40, 40
			        2574 => x"00000000",		-- colors: 40, 40, 40, 40
			        2575 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2576 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2577 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2578 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2579 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2580 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2581 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2582 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2583 => x"00000000",		-- colors: 40, 40, 40, 40
			        2584 => x"00000000",		-- colors: 40, 40, 40, 40
			        2585 => x"00000000",		-- colors: 40, 40, 40, 40
			        2586 => x"00000000",		-- colors: 40, 40, 40, 40
			        2587 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2588 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2589 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2590 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2591 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2592 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2593 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2594 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2595 => x"00000000",		-- colors: 40, 40, 40, 40
			        2596 => x"00000000",		-- colors: 40, 40, 40, 40
			        2597 => x"00000000",		-- colors: 40, 40, 40, 40
			        2598 => x"00000000",		-- colors: 40, 40, 40, 40
			        2599 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2600 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2601 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2602 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2603 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2604 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2605 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2606 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2607 => x"00000000",		-- colors: 40, 40, 40, 40
			        2608 => x"00000000",		-- colors: 40, 40, 40, 40
			        2609 => x"00000000",		-- colors: 40, 40, 40, 40
			        2610 => x"00000000",		-- colors: 40, 40, 40, 40
			        2611 => x"00000000",		-- colors: 40, 40, 40, 40
			        2612 => x"00000000",		-- colors: 40, 40, 40, 40
			        2613 => x"00000000",		-- colors: 40, 40, 40, 40
			        2614 => x"00000000",		-- colors: 40, 40, 40, 40
			        2615 => x"00000000",		-- colors: 40, 40, 40, 40
			        2616 => x"00000000",		-- colors: 40, 40, 40, 40
			        2617 => x"00000000",		-- colors: 40, 40, 40, 40
			        2618 => x"00000000",		-- colors: 40, 40, 40, 40
			        2619 => x"00000000",		-- colors: 40, 40, 40, 40
			        2620 => x"00000000",		-- colors: 40, 40, 40, 40
			        2621 => x"00000000",		-- colors: 40, 40, 40, 40
			        2622 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 37
			        2623 => x"00000000",		-- colors: 40, 40, 40, 40
			        2624 => x"00000000",		-- colors: 40, 40, 40, 40
			        2625 => x"00000000",		-- colors: 40, 40, 40, 40
			        2626 => x"00000000",		-- colors: 40, 40, 40, 40
			        2627 => x"00000000",		-- colors: 40, 40, 40, 40
			        2628 => x"00000000",		-- colors: 40, 40, 40, 40
			        2629 => x"00000000",		-- colors: 40, 40, 40, 40
			        2630 => x"00000000",		-- colors: 40, 40, 40, 40
			        2631 => x"00000000",		-- colors: 40, 40, 40, 40
			        2632 => x"00000000",		-- colors: 40, 40, 40, 40
			        2633 => x"00000000",		-- colors: 40, 40, 40, 40
			        2634 => x"00000000",		-- colors: 40, 40, 40, 40
			        2635 => x"00000000",		-- colors: 40, 40, 40, 40
			        2636 => x"00000000",		-- colors: 40, 40, 40, 40
			        2637 => x"00000000",		-- colors: 40, 40, 40, 40
			        2638 => x"00000000",		-- colors: 40, 40, 40, 40
			        2639 => x"00000000",		-- colors: 40, 40, 40, 40
			        2640 => x"00000000",		-- colors: 40, 40, 40, 40
			        2641 => x"00000000",		-- colors: 40, 40, 40, 40
			        2642 => x"00000000",		-- colors: 40, 40, 40, 40
			        2643 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2644 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2645 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2646 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2647 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2648 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2649 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2650 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2651 => x"00000000",		-- colors: 40, 40, 40, 40
			        2652 => x"00000000",		-- colors: 40, 40, 40, 40
			        2653 => x"00000000",		-- colors: 40, 40, 40, 40
			        2654 => x"00000000",		-- colors: 40, 40, 40, 40
			        2655 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2656 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2657 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2658 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2659 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2660 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2661 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2662 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2663 => x"00000000",		-- colors: 40, 40, 40, 40
			        2664 => x"00000000",		-- colors: 40, 40, 40, 40
			        2665 => x"00000000",		-- colors: 40, 40, 40, 40
			        2666 => x"00000000",		-- colors: 40, 40, 40, 40
			        2667 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2668 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2669 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2670 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2671 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2672 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2673 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2674 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2675 => x"00000000",		-- colors: 40, 40, 40, 40
			        2676 => x"00000000",		-- colors: 40, 40, 40, 40
			        2677 => x"00000000",		-- colors: 40, 40, 40, 40
			        2678 => x"00000000",		-- colors: 40, 40, 40, 40
			        2679 => x"32323232",		-- colors: 50, 50, 50, 50
			        2680 => x"32323232",		-- colors: 50, 50, 50, 50
			        2681 => x"32323232",		-- colors: 50, 50, 50, 50
			        2682 => x"32323232",		-- colors: 50, 50, 50, 50
			        2683 => x"00000000",		-- colors: 40, 40, 40, 40
			        2684 => x"00000000",		-- colors: 40, 40, 40, 40
			        2685 => x"00000000",		-- colors: 40, 40, 40, 40
			        2686 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 38
			        2687 => x"00000000",		-- colors: 40, 40, 40, 40
			        2688 => x"00000000",		-- colors: 40, 40, 40, 40
			        2689 => x"00000000",		-- colors: 40, 40, 40, 40
			        2690 => x"00000000",		-- colors: 40, 40, 40, 40
			        2691 => x"00000000",		-- colors: 40, 40, 40, 40
			        2692 => x"00000000",		-- colors: 40, 40, 40, 40
			        2693 => x"00000000",		-- colors: 40, 40, 40, 40
			        2694 => x"00000000",		-- colors: 40, 40, 40, 40
			        2695 => x"00000000",		-- colors: 40, 40, 40, 40
			        2696 => x"00000000",		-- colors: 40, 40, 40, 40
			        2697 => x"00000000",		-- colors: 40, 40, 40, 40
			        2698 => x"00000000",		-- colors: 40, 40, 40, 40
			        2699 => x"00000000",		-- colors: 40, 40, 40, 40
			        2700 => x"00000000",		-- colors: 40, 40, 40, 40
			        2701 => x"00000000",		-- colors: 40, 40, 40, 40
			        2702 => x"00000000",		-- colors: 40, 40, 40, 40
			        2703 => x"00000000",		-- colors: 40, 40, 40, 40
			        2704 => x"00000000",		-- colors: 40, 40, 40, 40
			        2705 => x"00000000",		-- colors: 40, 40, 40, 40
			        2706 => x"00000000",		-- colors: 40, 40, 40, 40
			        2707 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2708 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2709 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2710 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2711 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2712 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2713 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2714 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2715 => x"00000000",		-- colors: 40, 40, 40, 40
			        2716 => x"00000000",		-- colors: 40, 40, 40, 40
			        2717 => x"00000000",		-- colors: 40, 40, 40, 40
			        2718 => x"00000000",		-- colors: 40, 40, 40, 40
			        2719 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2720 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2721 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2722 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2723 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2724 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2725 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2726 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2727 => x"00000000",		-- colors: 40, 40, 40, 40
			        2728 => x"00000000",		-- colors: 40, 40, 40, 40
			        2729 => x"00000000",		-- colors: 40, 40, 40, 40
			        2730 => x"00000000",		-- colors: 40, 40, 40, 40
			        2731 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2732 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2733 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2734 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2735 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2736 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2737 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2738 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2739 => x"00000000",		-- colors: 40, 40, 40, 40
			        2740 => x"00000000",		-- colors: 40, 40, 40, 40
			        2741 => x"00000000",		-- colors: 40, 40, 40, 40
			        2742 => x"00000000",		-- colors: 40, 40, 40, 40
			        2743 => x"00000000",		-- colors: 40, 40, 40, 40
			        2744 => x"00000000",		-- colors: 40, 40, 40, 40
			        2745 => x"00000000",		-- colors: 40, 40, 40, 40
			        2746 => x"00000000",		-- colors: 40, 40, 40, 40
			        2747 => x"00000000",		-- colors: 40, 40, 40, 40
			        2748 => x"00000000",		-- colors: 40, 40, 40, 40
			        2749 => x"00000000",		-- colors: 40, 40, 40, 40
			        2750 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 39
			        2751 => x"00000000",		-- colors: 40, 40, 40, 40
			        2752 => x"00000000",		-- colors: 40, 40, 40, 40
			        2753 => x"00000000",		-- colors: 40, 40, 40, 40
			        2754 => x"00000000",		-- colors: 40, 40, 40, 40
			        2755 => x"00000000",		-- colors: 40, 40, 40, 40
			        2756 => x"00000000",		-- colors: 40, 40, 40, 40
			        2757 => x"00000000",		-- colors: 40, 40, 40, 40
			        2758 => x"00000000",		-- colors: 40, 40, 40, 40
			        2759 => x"00000000",		-- colors: 40, 40, 40, 40
			        2760 => x"00000000",		-- colors: 40, 40, 40, 40
			        2761 => x"00000000",		-- colors: 40, 40, 40, 40
			        2762 => x"00000000",		-- colors: 40, 40, 40, 40
			        2763 => x"00000000",		-- colors: 40, 40, 40, 40
			        2764 => x"00000000",		-- colors: 40, 40, 40, 40
			        2765 => x"00000000",		-- colors: 40, 40, 40, 40
			        2766 => x"00000000",		-- colors: 40, 40, 40, 40
			        2767 => x"00000000",		-- colors: 40, 40, 40, 40
			        2768 => x"00000000",		-- colors: 40, 40, 40, 40
			        2769 => x"00000000",		-- colors: 40, 40, 40, 40
			        2770 => x"00000000",		-- colors: 40, 40, 40, 40
			        2771 => x"00000000",		-- colors: 40, 40, 40, 40
			        2772 => x"00000000",		-- colors: 40, 40, 40, 40
			        2773 => x"00000000",		-- colors: 40, 40, 40, 40
			        2774 => x"00000000",		-- colors: 40, 40, 40, 40
			        2775 => x"00000000",		-- colors: 40, 40, 40, 40
			        2776 => x"00000000",		-- colors: 40, 40, 40, 40
			        2777 => x"00000000",		-- colors: 40, 40, 40, 40
			        2778 => x"00000000",		-- colors: 40, 40, 40, 40
			        2779 => x"00000000",		-- colors: 40, 40, 40, 40
			        2780 => x"00000000",		-- colors: 40, 40, 40, 40
			        2781 => x"00000000",		-- colors: 40, 40, 40, 40
			        2782 => x"00000000",		-- colors: 40, 40, 40, 40
			        2783 => x"00000000",		-- colors: 40, 40, 40, 40
			        2784 => x"00000000",		-- colors: 40, 40, 40, 40
			        2785 => x"00000000",		-- colors: 40, 40, 40, 40
			        2786 => x"00000000",		-- colors: 40, 40, 40, 40
			        2787 => x"00000000",		-- colors: 40, 40, 40, 40
			        2788 => x"00000000",		-- colors: 40, 40, 40, 40
			        2789 => x"00000000",		-- colors: 40, 40, 40, 40
			        2790 => x"00000000",		-- colors: 40, 40, 40, 40
			        2791 => x"32323232",		-- colors: 50, 50, 50, 50
			        2792 => x"32323232",		-- colors: 50, 50, 50, 50
			        2793 => x"32323232",		-- colors: 50, 50, 50, 50
			        2794 => x"32323232",		-- colors: 50, 50, 50, 50
			        2795 => x"00000000",		-- colors: 40, 40, 40, 40
			        2796 => x"00000000",		-- colors: 40, 40, 40, 40
			        2797 => x"00000000",		-- colors: 40, 40, 40, 40
			        2798 => x"00000000",		-- colors: 40, 40, 40, 40
			        2799 => x"00000000",		-- colors: 40, 40, 40, 40
			        2800 => x"00000000",		-- colors: 40, 40, 40, 40
			        2801 => x"00000000",		-- colors: 40, 40, 40, 40
			        2802 => x"00000000",		-- colors: 40, 40, 40, 40
			        2803 => x"00000000",		-- colors: 40, 40, 40, 40
			        2804 => x"00000000",		-- colors: 40, 40, 40, 40
			        2805 => x"00000000",		-- colors: 40, 40, 40, 40
			        2806 => x"00000000",		-- colors: 40, 40, 40, 40
			        2807 => x"32323232",		-- colors: 50, 50, 50, 50
			        2808 => x"32323232",		-- colors: 50, 50, 50, 50
			        2809 => x"32323232",		-- colors: 50, 50, 50, 50
			        2810 => x"32323232",		-- colors: 50, 50, 50, 50
			        2811 => x"00000000",		-- colors: 40, 40, 40, 40
			        2812 => x"00000000",		-- colors: 40, 40, 40, 40
			        2813 => x"00000000",		-- colors: 40, 40, 40, 40
			        2814 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 40
			        2815 => x"00000000",		-- colors: 40, 40, 40, 40
			        2816 => x"00000000",		-- colors: 40, 40, 40, 40
			        2817 => x"00000000",		-- colors: 40, 40, 40, 40
			        2818 => x"00000000",		-- colors: 40, 40, 40, 40
			        2819 => x"00000000",		-- colors: 40, 40, 40, 40
			        2820 => x"00000000",		-- colors: 40, 40, 40, 40
			        2821 => x"00000000",		-- colors: 40, 40, 40, 40
			        2822 => x"00000000",		-- colors: 40, 40, 40, 40
			        2823 => x"00000000",		-- colors: 40, 40, 40, 40
			        2824 => x"00000000",		-- colors: 40, 40, 40, 40
			        2825 => x"00000000",		-- colors: 40, 40, 40, 40
			        2826 => x"00000000",		-- colors: 40, 40, 40, 40
			        2827 => x"00000000",		-- colors: 40, 40, 40, 40
			        2828 => x"00000000",		-- colors: 40, 40, 40, 40
			        2829 => x"00000000",		-- colors: 40, 40, 40, 40
			        2830 => x"00000000",		-- colors: 40, 40, 40, 40
			        2831 => x"00000000",		-- colors: 40, 40, 40, 40
			        2832 => x"00000000",		-- colors: 40, 40, 40, 40
			        2833 => x"00000000",		-- colors: 40, 40, 40, 40
			        2834 => x"00000000",		-- colors: 40, 40, 40, 40
			        2835 => x"00000000",		-- colors: 40, 40, 40, 40
			        2836 => x"00000000",		-- colors: 40, 40, 40, 40
			        2837 => x"00000000",		-- colors: 40, 40, 40, 40
			        2838 => x"00000000",		-- colors: 40, 40, 40, 40
			        2839 => x"00000000",		-- colors: 40, 40, 40, 40
			        2840 => x"00000000",		-- colors: 40, 40, 40, 40
			        2841 => x"00000000",		-- colors: 40, 40, 40, 40
			        2842 => x"00000000",		-- colors: 40, 40, 40, 40
			        2843 => x"00000000",		-- colors: 40, 40, 40, 40
			        2844 => x"00000000",		-- colors: 40, 40, 40, 40
			        2845 => x"00000000",		-- colors: 40, 40, 40, 40
			        2846 => x"00000000",		-- colors: 40, 40, 40, 40
			        2847 => x"00000000",		-- colors: 40, 40, 40, 40
			        2848 => x"00000000",		-- colors: 40, 40, 40, 40
			        2849 => x"00000000",		-- colors: 40, 40, 40, 40
			        2850 => x"00000000",		-- colors: 40, 40, 40, 40
			        2851 => x"00000000",		-- colors: 40, 40, 40, 40
			        2852 => x"00000000",		-- colors: 40, 40, 40, 40
			        2853 => x"00000000",		-- colors: 40, 40, 40, 40
			        2854 => x"00000000",		-- colors: 40, 40, 40, 40
			        2855 => x"00000000",		-- colors: 40, 40, 40, 40
			        2856 => x"00000000",		-- colors: 40, 40, 40, 40
			        2857 => x"00000000",		-- colors: 40, 40, 40, 40
			        2858 => x"00000000",		-- colors: 40, 40, 40, 40
			        2859 => x"00000000",		-- colors: 40, 40, 40, 40
			        2860 => x"00000000",		-- colors: 40, 40, 40, 40
			        2861 => x"00000000",		-- colors: 40, 40, 40, 40
			        2862 => x"00000000",		-- colors: 40, 40, 40, 40
			        2863 => x"00000000",		-- colors: 40, 40, 40, 40
			        2864 => x"00000000",		-- colors: 40, 40, 40, 40
			        2865 => x"00000000",		-- colors: 40, 40, 40, 40
			        2866 => x"00000000",		-- colors: 40, 40, 40, 40
			        2867 => x"00000000",		-- colors: 40, 40, 40, 40
			        2868 => x"00000000",		-- colors: 40, 40, 40, 40
			        2869 => x"00000000",		-- colors: 40, 40, 40, 40
			        2870 => x"00000000",		-- colors: 40, 40, 40, 40
			        2871 => x"00000000",		-- colors: 40, 40, 40, 40
			        2872 => x"00000000",		-- colors: 40, 40, 40, 40
			        2873 => x"00000000",		-- colors: 40, 40, 40, 40
			        2874 => x"00000000",		-- colors: 40, 40, 40, 40
			        2875 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2876 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2877 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2878 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60

			                --  sprite 41
			        2879 => x"00000000",		-- colors: 40, 40, 40, 40
			        2880 => x"00000000",		-- colors: 40, 40, 40, 40
			        2881 => x"00000000",		-- colors: 40, 40, 40, 40
			        2882 => x"00000000",		-- colors: 40, 40, 40, 40
			        2883 => x"00000000",		-- colors: 40, 40, 40, 40
			        2884 => x"00000000",		-- colors: 40, 40, 40, 40
			        2885 => x"00000000",		-- colors: 40, 40, 40, 40
			        2886 => x"00000000",		-- colors: 40, 40, 40, 40
			        2887 => x"00000000",		-- colors: 40, 40, 40, 40
			        2888 => x"00000000",		-- colors: 40, 40, 40, 40
			        2889 => x"00000000",		-- colors: 40, 40, 40, 40
			        2890 => x"00000000",		-- colors: 40, 40, 40, 40
			        2891 => x"00000000",		-- colors: 40, 40, 40, 40
			        2892 => x"00000000",		-- colors: 40, 40, 40, 40
			        2893 => x"00000000",		-- colors: 40, 40, 40, 40
			        2894 => x"00000000",		-- colors: 40, 40, 40, 40
			        2895 => x"00000000",		-- colors: 40, 40, 40, 40
			        2896 => x"00000000",		-- colors: 40, 40, 40, 40
			        2897 => x"00000000",		-- colors: 40, 40, 40, 40
			        2898 => x"00000000",		-- colors: 40, 40, 40, 40
			        2899 => x"00000000",		-- colors: 40, 40, 40, 40
			        2900 => x"00000000",		-- colors: 40, 40, 40, 40
			        2901 => x"00000000",		-- colors: 40, 40, 40, 40
			        2902 => x"00000000",		-- colors: 40, 40, 40, 40
			        2903 => x"00000000",		-- colors: 40, 40, 40, 40
			        2904 => x"00000000",		-- colors: 40, 40, 40, 40
			        2905 => x"00000000",		-- colors: 40, 40, 40, 40
			        2906 => x"00000000",		-- colors: 40, 40, 40, 40
			        2907 => x"00000000",		-- colors: 40, 40, 40, 40
			        2908 => x"00000000",		-- colors: 40, 40, 40, 40
			        2909 => x"00000000",		-- colors: 40, 40, 40, 40
			        2910 => x"00000000",		-- colors: 40, 40, 40, 40
			        2911 => x"00000000",		-- colors: 40, 40, 40, 40
			        2912 => x"00000000",		-- colors: 40, 40, 40, 40
			        2913 => x"00000000",		-- colors: 40, 40, 40, 40
			        2914 => x"00000000",		-- colors: 40, 40, 40, 40
			        2915 => x"00000000",		-- colors: 40, 40, 40, 40
			        2916 => x"00000000",		-- colors: 40, 40, 40, 40
			        2917 => x"00000000",		-- colors: 40, 40, 40, 40
			        2918 => x"00000000",		-- colors: 40, 40, 40, 40
			        2919 => x"00000000",		-- colors: 40, 40, 40, 40
			        2920 => x"00000000",		-- colors: 40, 40, 40, 40
			        2921 => x"00000000",		-- colors: 40, 40, 40, 40
			        2922 => x"00000000",		-- colors: 40, 40, 40, 40
			        2923 => x"00000000",		-- colors: 40, 40, 40, 40
			        2924 => x"00000000",		-- colors: 40, 40, 40, 40
			        2925 => x"00000000",		-- colors: 40, 40, 40, 40
			        2926 => x"00000000",		-- colors: 40, 40, 40, 40
			        2927 => x"00000000",		-- colors: 40, 40, 40, 40
			        2928 => x"00000000",		-- colors: 40, 40, 40, 40
			        2929 => x"00000000",		-- colors: 40, 40, 40, 40
			        2930 => x"00000000",		-- colors: 40, 40, 40, 40
			        2931 => x"00000000",		-- colors: 40, 40, 40, 40
			        2932 => x"00000000",		-- colors: 40, 40, 40, 40
			        2933 => x"00000000",		-- colors: 40, 40, 40, 40
			        2934 => x"00000000",		-- colors: 40, 40, 40, 40
			        2935 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2936 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2937 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2938 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2939 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2940 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2941 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        2942 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60

			                --  sprite 42
			        2943 => x"00000000",		-- colors: 40, 40, 40, 40
			        2944 => x"00000000",		-- colors: 40, 40, 40, 40
			        2945 => x"00000000",		-- colors: 40, 40, 40, 40
			        2946 => x"00000000",		-- colors: 40, 40, 40, 40
			        2947 => x"00000000",		-- colors: 40, 40, 40, 40
			        2948 => x"00000000",		-- colors: 40, 40, 40, 40
			        2949 => x"00000000",		-- colors: 40, 40, 40, 40
			        2950 => x"00000000",		-- colors: 40, 40, 40, 40
			        2951 => x"00000000",		-- colors: 40, 40, 40, 40
			        2952 => x"00000000",		-- colors: 40, 40, 40, 40
			        2953 => x"00000000",		-- colors: 40, 40, 40, 40
			        2954 => x"00000000",		-- colors: 40, 40, 40, 40
			        2955 => x"00000000",		-- colors: 40, 40, 40, 40
			        2956 => x"00000000",		-- colors: 40, 40, 40, 40
			        2957 => x"00000000",		-- colors: 40, 40, 40, 40
			        2958 => x"00000000",		-- colors: 40, 40, 40, 40
			        2959 => x"00000000",		-- colors: 40, 40, 40, 40
			        2960 => x"00000000",		-- colors: 40, 40, 40, 40
			        2961 => x"00000000",		-- colors: 40, 40, 40, 40
			        2962 => x"00000000",		-- colors: 40, 40, 40, 40
			        2963 => x"00000000",		-- colors: 40, 40, 40, 40
			        2964 => x"00000000",		-- colors: 40, 40, 40, 40
			        2965 => x"00000000",		-- colors: 40, 40, 40, 40
			        2966 => x"00000000",		-- colors: 40, 40, 40, 40
			        2967 => x"00000000",		-- colors: 40, 40, 40, 40
			        2968 => x"00000000",		-- colors: 40, 40, 40, 40
			        2969 => x"00000000",		-- colors: 40, 40, 40, 40
			        2970 => x"00000000",		-- colors: 40, 40, 40, 40
			        2971 => x"00000000",		-- colors: 40, 40, 40, 40
			        2972 => x"00000000",		-- colors: 40, 40, 40, 40
			        2973 => x"00000000",		-- colors: 40, 40, 40, 40
			        2974 => x"00000000",		-- colors: 40, 40, 40, 40
			        2975 => x"00000000",		-- colors: 40, 40, 40, 40
			        2976 => x"00000000",		-- colors: 40, 40, 40, 40
			        2977 => x"00000000",		-- colors: 40, 40, 40, 40
			        2978 => x"00000000",		-- colors: 40, 40, 40, 40
			        2979 => x"00000000",		-- colors: 40, 40, 40, 40
			        2980 => x"00000000",		-- colors: 40, 40, 40, 40
			        2981 => x"00000000",		-- colors: 40, 40, 40, 40
			        2982 => x"00000000",		-- colors: 40, 40, 40, 40
			        2983 => x"00000000",		-- colors: 40, 40, 40, 40
			        2984 => x"00000000",		-- colors: 40, 40, 40, 40
			        2985 => x"00000000",		-- colors: 40, 40, 40, 40
			        2986 => x"00000000",		-- colors: 40, 40, 40, 40
			        2987 => x"00000000",		-- colors: 40, 40, 40, 40
			        2988 => x"00000000",		-- colors: 40, 40, 40, 40
			        2989 => x"00000000",		-- colors: 40, 40, 40, 40
			        2990 => x"00000000",		-- colors: 40, 40, 40, 40
			        2991 => x"00000000",		-- colors: 40, 40, 40, 40
			        2992 => x"00000000",		-- colors: 40, 40, 40, 40
			        2993 => x"00000000",		-- colors: 40, 40, 40, 40
			        2994 => x"00000000",		-- colors: 40, 40, 40, 40
			        2995 => x"00000000",		-- colors: 40, 40, 40, 40
			        2996 => x"00000000",		-- colors: 40, 40, 40, 40
			        2997 => x"00000000",		-- colors: 40, 40, 40, 40
			        2998 => x"00000000",		-- colors: 40, 40, 40, 40
			        2999 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3000 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3001 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3002 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3003 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3004 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3005 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3006 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60

			                --  sprite 43
			        3007 => x"00000000",		-- colors: 40, 40, 40, 40
			        3008 => x"00000000",		-- colors: 40, 40, 40, 40
			        3009 => x"00000000",		-- colors: 40, 40, 40, 40
			        3010 => x"00000000",		-- colors: 40, 40, 40, 40
			        3011 => x"00000000",		-- colors: 40, 40, 40, 40
			        3012 => x"00000000",		-- colors: 40, 40, 40, 40
			        3013 => x"00000000",		-- colors: 40, 40, 40, 40
			        3014 => x"00000000",		-- colors: 40, 40, 40, 40
			        3015 => x"00000000",		-- colors: 40, 40, 40, 40
			        3016 => x"00000000",		-- colors: 40, 40, 40, 40
			        3017 => x"00000000",		-- colors: 40, 40, 40, 40
			        3018 => x"00000000",		-- colors: 40, 40, 40, 40
			        3019 => x"00000000",		-- colors: 40, 40, 40, 40
			        3020 => x"00000000",		-- colors: 40, 40, 40, 40
			        3021 => x"00000000",		-- colors: 40, 40, 40, 40
			        3022 => x"00000000",		-- colors: 40, 40, 40, 40
			        3023 => x"00000000",		-- colors: 40, 40, 40, 40
			        3024 => x"00000000",		-- colors: 40, 40, 40, 40
			        3025 => x"00000000",		-- colors: 40, 40, 40, 40
			        3026 => x"00000000",		-- colors: 40, 40, 40, 40
			        3027 => x"00000000",		-- colors: 40, 40, 40, 40
			        3028 => x"00000000",		-- colors: 40, 40, 40, 40
			        3029 => x"00000000",		-- colors: 40, 40, 40, 40
			        3030 => x"00000000",		-- colors: 40, 40, 40, 40
			        3031 => x"00000000",		-- colors: 40, 40, 40, 40
			        3032 => x"00000000",		-- colors: 40, 40, 40, 40
			        3033 => x"00000000",		-- colors: 40, 40, 40, 40
			        3034 => x"00000000",		-- colors: 40, 40, 40, 40
			        3035 => x"00000000",		-- colors: 40, 40, 40, 40
			        3036 => x"00000000",		-- colors: 40, 40, 40, 40
			        3037 => x"00000000",		-- colors: 40, 40, 40, 40
			        3038 => x"00000000",		-- colors: 40, 40, 40, 40
			        3039 => x"00000000",		-- colors: 40, 40, 40, 40
			        3040 => x"00000000",		-- colors: 40, 40, 40, 40
			        3041 => x"00000000",		-- colors: 40, 40, 40, 40
			        3042 => x"00000000",		-- colors: 40, 40, 40, 40
			        3043 => x"00000000",		-- colors: 40, 40, 40, 40
			        3044 => x"00000000",		-- colors: 40, 40, 40, 40
			        3045 => x"00000000",		-- colors: 40, 40, 40, 40
			        3046 => x"00000000",		-- colors: 40, 40, 40, 40
			        3047 => x"00000000",		-- colors: 40, 40, 40, 40
			        3048 => x"00000000",		-- colors: 40, 40, 40, 40
			        3049 => x"00000000",		-- colors: 40, 40, 40, 40
			        3050 => x"00000000",		-- colors: 40, 40, 40, 40
			        3051 => x"00000000",		-- colors: 40, 40, 40, 40
			        3052 => x"00000000",		-- colors: 40, 40, 40, 40
			        3053 => x"00000000",		-- colors: 40, 40, 40, 40
			        3054 => x"00000000",		-- colors: 40, 40, 40, 40
			        3055 => x"00000000",		-- colors: 40, 40, 40, 40
			        3056 => x"00000000",		-- colors: 40, 40, 40, 40
			        3057 => x"00000000",		-- colors: 40, 40, 40, 40
			        3058 => x"00000000",		-- colors: 40, 40, 40, 40
			        3059 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3060 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3061 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3062 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3063 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3064 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3065 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3066 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3067 => x"00000000",		-- colors: 40, 40, 40, 40
			        3068 => x"00000000",		-- colors: 40, 40, 40, 40
			        3069 => x"00000000",		-- colors: 40, 40, 40, 40
			        3070 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 44
			        3071 => x"00000000",		-- colors: 40, 40, 40, 40
			        3072 => x"00000000",		-- colors: 40, 40, 40, 40
			        3073 => x"00000000",		-- colors: 40, 40, 40, 40
			        3074 => x"00000000",		-- colors: 40, 40, 40, 40
			        3075 => x"00000000",		-- colors: 40, 40, 40, 40
			        3076 => x"00000000",		-- colors: 40, 40, 40, 40
			        3077 => x"00000000",		-- colors: 40, 40, 40, 40
			        3078 => x"00000000",		-- colors: 40, 40, 40, 40
			        3079 => x"32323232",		-- colors: 50, 50, 50, 50
			        3080 => x"32323232",		-- colors: 50, 50, 50, 50
			        3081 => x"32323232",		-- colors: 50, 50, 50, 50
			        3082 => x"32323232",		-- colors: 50, 50, 50, 50
			        3083 => x"00000000",		-- colors: 40, 40, 40, 40
			        3084 => x"00000000",		-- colors: 40, 40, 40, 40
			        3085 => x"00000000",		-- colors: 40, 40, 40, 40
			        3086 => x"00000000",		-- colors: 40, 40, 40, 40
			        3087 => x"00000000",		-- colors: 40, 40, 40, 40
			        3088 => x"00000000",		-- colors: 40, 40, 40, 40
			        3089 => x"00000000",		-- colors: 40, 40, 40, 40
			        3090 => x"00000000",		-- colors: 40, 40, 40, 40
			        3091 => x"00000000",		-- colors: 40, 40, 40, 40
			        3092 => x"00000000",		-- colors: 40, 40, 40, 40
			        3093 => x"00000000",		-- colors: 40, 40, 40, 40
			        3094 => x"00000000",		-- colors: 40, 40, 40, 40
			        3095 => x"32323232",		-- colors: 50, 50, 50, 50
			        3096 => x"32323232",		-- colors: 50, 50, 50, 50
			        3097 => x"32323232",		-- colors: 50, 50, 50, 50
			        3098 => x"32323232",		-- colors: 50, 50, 50, 50
			        3099 => x"00000000",		-- colors: 40, 40, 40, 40
			        3100 => x"00000000",		-- colors: 40, 40, 40, 40
			        3101 => x"00000000",		-- colors: 40, 40, 40, 40
			        3102 => x"00000000",		-- colors: 40, 40, 40, 40
			        3103 => x"00000000",		-- colors: 40, 40, 40, 40
			        3104 => x"00000000",		-- colors: 40, 40, 40, 40
			        3105 => x"00000000",		-- colors: 40, 40, 40, 40
			        3106 => x"00000000",		-- colors: 40, 40, 40, 40
			        3107 => x"00000000",		-- colors: 40, 40, 40, 40
			        3108 => x"00000000",		-- colors: 40, 40, 40, 40
			        3109 => x"00000000",		-- colors: 40, 40, 40, 40
			        3110 => x"00000000",		-- colors: 40, 40, 40, 40
			        3111 => x"32323232",		-- colors: 50, 50, 50, 50
			        3112 => x"32323232",		-- colors: 50, 50, 50, 50
			        3113 => x"32323232",		-- colors: 50, 50, 50, 50
			        3114 => x"32323232",		-- colors: 50, 50, 50, 50
			        3115 => x"00000000",		-- colors: 40, 40, 40, 40
			        3116 => x"00000000",		-- colors: 40, 40, 40, 40
			        3117 => x"00000000",		-- colors: 40, 40, 40, 40
			        3118 => x"00000000",		-- colors: 40, 40, 40, 40
			        3119 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3120 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3121 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3122 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3123 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3124 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3125 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3126 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3127 => x"00000000",		-- colors: 40, 40, 40, 40
			        3128 => x"00000000",		-- colors: 40, 40, 40, 40
			        3129 => x"00000000",		-- colors: 40, 40, 40, 40
			        3130 => x"00000000",		-- colors: 40, 40, 40, 40
			        3131 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3132 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3133 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3134 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60

			                --  sprite 45
			        3135 => x"00000000",		-- colors: 40, 40, 40, 40
			        3136 => x"00000000",		-- colors: 40, 40, 40, 40
			        3137 => x"00000000",		-- colors: 40, 40, 40, 40
			        3138 => x"00000000",		-- colors: 40, 40, 40, 40
			        3139 => x"00000000",		-- colors: 40, 40, 40, 40
			        3140 => x"00000000",		-- colors: 40, 40, 40, 40
			        3141 => x"00000000",		-- colors: 40, 40, 40, 40
			        3142 => x"00000000",		-- colors: 40, 40, 40, 40
			        3143 => x"00000000",		-- colors: 40, 40, 40, 40
			        3144 => x"00000000",		-- colors: 40, 40, 40, 40
			        3145 => x"00000000",		-- colors: 40, 40, 40, 40
			        3146 => x"00000000",		-- colors: 40, 40, 40, 40
			        3147 => x"00000000",		-- colors: 40, 40, 40, 40
			        3148 => x"00000000",		-- colors: 40, 40, 40, 40
			        3149 => x"00000000",		-- colors: 40, 40, 40, 40
			        3150 => x"00000000",		-- colors: 40, 40, 40, 40
			        3151 => x"00000000",		-- colors: 40, 40, 40, 40
			        3152 => x"00000000",		-- colors: 40, 40, 40, 40
			        3153 => x"00000000",		-- colors: 40, 40, 40, 40
			        3154 => x"00000000",		-- colors: 40, 40, 40, 40
			        3155 => x"00000000",		-- colors: 40, 40, 40, 40
			        3156 => x"00000000",		-- colors: 40, 40, 40, 40
			        3157 => x"00000000",		-- colors: 40, 40, 40, 40
			        3158 => x"00000000",		-- colors: 40, 40, 40, 40
			        3159 => x"00000000",		-- colors: 40, 40, 40, 40
			        3160 => x"00000000",		-- colors: 40, 40, 40, 40
			        3161 => x"00000000",		-- colors: 40, 40, 40, 40
			        3162 => x"00000000",		-- colors: 40, 40, 40, 40
			        3163 => x"00000000",		-- colors: 40, 40, 40, 40
			        3164 => x"00000000",		-- colors: 40, 40, 40, 40
			        3165 => x"00000000",		-- colors: 40, 40, 40, 40
			        3166 => x"00000000",		-- colors: 40, 40, 40, 40
			        3167 => x"00000000",		-- colors: 40, 40, 40, 40
			        3168 => x"00000000",		-- colors: 40, 40, 40, 40
			        3169 => x"00000000",		-- colors: 40, 40, 40, 40
			        3170 => x"00000000",		-- colors: 40, 40, 40, 40
			        3171 => x"00000000",		-- colors: 40, 40, 40, 40
			        3172 => x"00000000",		-- colors: 40, 40, 40, 40
			        3173 => x"00000000",		-- colors: 40, 40, 40, 40
			        3174 => x"00000000",		-- colors: 40, 40, 40, 40
			        3175 => x"00000000",		-- colors: 40, 40, 40, 40
			        3176 => x"00000000",		-- colors: 40, 40, 40, 40
			        3177 => x"00000000",		-- colors: 40, 40, 40, 40
			        3178 => x"00000000",		-- colors: 40, 40, 40, 40
			        3179 => x"00000000",		-- colors: 40, 40, 40, 40
			        3180 => x"00000000",		-- colors: 40, 40, 40, 40
			        3181 => x"00000000",		-- colors: 40, 40, 40, 40
			        3182 => x"00000000",		-- colors: 40, 40, 40, 40
			        3183 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3184 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3185 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3186 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3187 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3188 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3189 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3190 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3191 => x"00000000",		-- colors: 40, 40, 40, 40
			        3192 => x"00000000",		-- colors: 40, 40, 40, 40
			        3193 => x"00000000",		-- colors: 40, 40, 40, 40
			        3194 => x"00000000",		-- colors: 40, 40, 40, 40
			        3195 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3196 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3197 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3198 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60

			                --  sprite 46
			        3199 => x"00000000",		-- colors: 40, 40, 40, 40
			        3200 => x"00000000",		-- colors: 40, 40, 40, 40
			        3201 => x"00000000",		-- colors: 40, 40, 40, 40
			        3202 => x"00000000",		-- colors: 40, 40, 40, 40
			        3203 => x"00000000",		-- colors: 40, 40, 40, 40
			        3204 => x"00000000",		-- colors: 40, 40, 40, 40
			        3205 => x"00000000",		-- colors: 40, 40, 40, 40
			        3206 => x"00000000",		-- colors: 40, 40, 40, 40
			        3207 => x"00000000",		-- colors: 40, 40, 40, 40
			        3208 => x"00000000",		-- colors: 40, 40, 40, 40
			        3209 => x"00000000",		-- colors: 40, 40, 40, 40
			        3210 => x"00000000",		-- colors: 40, 40, 40, 40
			        3211 => x"00000000",		-- colors: 40, 40, 40, 40
			        3212 => x"00000000",		-- colors: 40, 40, 40, 40
			        3213 => x"00000000",		-- colors: 40, 40, 40, 40
			        3214 => x"00000000",		-- colors: 40, 40, 40, 40
			        3215 => x"00000000",		-- colors: 40, 40, 40, 40
			        3216 => x"00000000",		-- colors: 40, 40, 40, 40
			        3217 => x"00000000",		-- colors: 40, 40, 40, 40
			        3218 => x"00000000",		-- colors: 40, 40, 40, 40
			        3219 => x"00000000",		-- colors: 40, 40, 40, 40
			        3220 => x"00000000",		-- colors: 40, 40, 40, 40
			        3221 => x"00000000",		-- colors: 40, 40, 40, 40
			        3222 => x"00000000",		-- colors: 40, 40, 40, 40
			        3223 => x"00000000",		-- colors: 40, 40, 40, 40
			        3224 => x"00000000",		-- colors: 40, 40, 40, 40
			        3225 => x"00000000",		-- colors: 40, 40, 40, 40
			        3226 => x"00000000",		-- colors: 40, 40, 40, 40
			        3227 => x"00000000",		-- colors: 40, 40, 40, 40
			        3228 => x"00000000",		-- colors: 40, 40, 40, 40
			        3229 => x"00000000",		-- colors: 40, 40, 40, 40
			        3230 => x"00000000",		-- colors: 40, 40, 40, 40
			        3231 => x"00000000",		-- colors: 40, 40, 40, 40
			        3232 => x"00000000",		-- colors: 40, 40, 40, 40
			        3233 => x"00000000",		-- colors: 40, 40, 40, 40
			        3234 => x"00000000",		-- colors: 40, 40, 40, 40
			        3235 => x"00000000",		-- colors: 40, 40, 40, 40
			        3236 => x"00000000",		-- colors: 40, 40, 40, 40
			        3237 => x"00000000",		-- colors: 40, 40, 40, 40
			        3238 => x"00000000",		-- colors: 40, 40, 40, 40
			        3239 => x"00000000",		-- colors: 40, 40, 40, 40
			        3240 => x"00000000",		-- colors: 40, 40, 40, 40
			        3241 => x"00000000",		-- colors: 40, 40, 40, 40
			        3242 => x"00000000",		-- colors: 40, 40, 40, 40
			        3243 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3244 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3245 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3246 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3247 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3248 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3249 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3250 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3251 => x"00000000",		-- colors: 40, 40, 40, 40
			        3252 => x"00000000",		-- colors: 40, 40, 40, 40
			        3253 => x"00000000",		-- colors: 40, 40, 40, 40
			        3254 => x"00000000",		-- colors: 40, 40, 40, 40
			        3255 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3256 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3257 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3258 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3259 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3260 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3261 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3262 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60

			                --  sprite 47
			        3263 => x"00000000",		-- colors: 40, 40, 40, 40
			        3264 => x"00000000",		-- colors: 40, 40, 40, 40
			        3265 => x"00000000",		-- colors: 40, 40, 40, 40
			        3266 => x"00000000",		-- colors: 40, 40, 40, 40
			        3267 => x"00000000",		-- colors: 40, 40, 40, 40
			        3268 => x"00000000",		-- colors: 40, 40, 40, 40
			        3269 => x"00000000",		-- colors: 40, 40, 40, 40
			        3270 => x"00000000",		-- colors: 40, 40, 40, 40
			        3271 => x"00000000",		-- colors: 40, 40, 40, 40
			        3272 => x"00000000",		-- colors: 40, 40, 40, 40
			        3273 => x"00000000",		-- colors: 40, 40, 40, 40
			        3274 => x"00000000",		-- colors: 40, 40, 40, 40
			        3275 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3276 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3277 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3278 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3279 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3280 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3281 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3282 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3283 => x"00000000",		-- colors: 40, 40, 40, 40
			        3284 => x"00000000",		-- colors: 40, 40, 40, 40
			        3285 => x"00000000",		-- colors: 40, 40, 40, 40
			        3286 => x"00000000",		-- colors: 40, 40, 40, 40
			        3287 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3288 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3289 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3290 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3291 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3292 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3293 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3294 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3295 => x"00000000",		-- colors: 40, 40, 40, 40
			        3296 => x"00000000",		-- colors: 40, 40, 40, 40
			        3297 => x"00000000",		-- colors: 40, 40, 40, 40
			        3298 => x"00000000",		-- colors: 40, 40, 40, 40
			        3299 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3300 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3301 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3302 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3303 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3304 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3305 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3306 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3307 => x"00000000",		-- colors: 40, 40, 40, 40
			        3308 => x"00000000",		-- colors: 40, 40, 40, 40
			        3309 => x"00000000",		-- colors: 40, 40, 40, 40
			        3310 => x"00000000",		-- colors: 40, 40, 40, 40
			        3311 => x"00000000",		-- colors: 40, 40, 40, 40
			        3312 => x"00000000",		-- colors: 40, 40, 40, 40
			        3313 => x"00000000",		-- colors: 40, 40, 40, 40
			        3314 => x"00000000",		-- colors: 40, 40, 40, 40
			        3315 => x"00000000",		-- colors: 40, 40, 40, 40
			        3316 => x"00000000",		-- colors: 40, 40, 40, 40
			        3317 => x"00000000",		-- colors: 40, 40, 40, 40
			        3318 => x"00000000",		-- colors: 40, 40, 40, 40
			        3319 => x"00000000",		-- colors: 40, 40, 40, 40
			        3320 => x"00000000",		-- colors: 40, 40, 40, 40
			        3321 => x"00000000",		-- colors: 40, 40, 40, 40
			        3322 => x"00000000",		-- colors: 40, 40, 40, 40
			        3323 => x"00000000",		-- colors: 40, 40, 40, 40
			        3324 => x"00000000",		-- colors: 40, 40, 40, 40
			        3325 => x"00000000",		-- colors: 40, 40, 40, 40
			        3326 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 48
			        3327 => x"00000000",		-- colors: 40, 40, 40, 40
			        3328 => x"00000000",		-- colors: 40, 40, 40, 40
			        3329 => x"00000000",		-- colors: 40, 40, 40, 40
			        3330 => x"00000000",		-- colors: 40, 40, 40, 40
			        3331 => x"00000000",		-- colors: 40, 40, 40, 40
			        3332 => x"00000000",		-- colors: 40, 40, 40, 40
			        3333 => x"00000000",		-- colors: 40, 40, 40, 40
			        3334 => x"00000000",		-- colors: 40, 40, 40, 40
			        3335 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3336 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3337 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3338 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3339 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3340 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3341 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3342 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3343 => x"00000000",		-- colors: 40, 40, 40, 40
			        3344 => x"00000000",		-- colors: 40, 40, 40, 40
			        3345 => x"00000000",		-- colors: 40, 40, 40, 40
			        3346 => x"00000000",		-- colors: 40, 40, 40, 40
			        3347 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3348 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3349 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3350 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3351 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3352 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3353 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3354 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3355 => x"00000000",		-- colors: 40, 40, 40, 40
			        3356 => x"00000000",		-- colors: 40, 40, 40, 40
			        3357 => x"00000000",		-- colors: 40, 40, 40, 40
			        3358 => x"00000000",		-- colors: 40, 40, 40, 40
			        3359 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3360 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3361 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3362 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3363 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3364 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3365 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3366 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3367 => x"00000000",		-- colors: 40, 40, 40, 40
			        3368 => x"00000000",		-- colors: 40, 40, 40, 40
			        3369 => x"00000000",		-- colors: 40, 40, 40, 40
			        3370 => x"00000000",		-- colors: 40, 40, 40, 40
			        3371 => x"00000000",		-- colors: 40, 40, 40, 40
			        3372 => x"00000000",		-- colors: 40, 40, 40, 40
			        3373 => x"00000000",		-- colors: 40, 40, 40, 40
			        3374 => x"00000000",		-- colors: 40, 40, 40, 40
			        3375 => x"00000000",		-- colors: 40, 40, 40, 40
			        3376 => x"00000000",		-- colors: 40, 40, 40, 40
			        3377 => x"00000000",		-- colors: 40, 40, 40, 40
			        3378 => x"00000000",		-- colors: 40, 40, 40, 40
			        3379 => x"00000000",		-- colors: 40, 40, 40, 40
			        3380 => x"00000000",		-- colors: 40, 40, 40, 40
			        3381 => x"00000000",		-- colors: 40, 40, 40, 40
			        3382 => x"00000000",		-- colors: 40, 40, 40, 40
			        3383 => x"00000000",		-- colors: 40, 40, 40, 40
			        3384 => x"00000000",		-- colors: 40, 40, 40, 40
			        3385 => x"00000000",		-- colors: 40, 40, 40, 40
			        3386 => x"00000000",		-- colors: 40, 40, 40, 40
			        3387 => x"00000000",		-- colors: 40, 40, 40, 40
			        3388 => x"00000000",		-- colors: 40, 40, 40, 40
			        3389 => x"00000000",		-- colors: 40, 40, 40, 40
			        3390 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 49
			        3391 => x"00000000",		-- colors: 40, 40, 40, 40
			        3392 => x"00000000",		-- colors: 40, 40, 40, 40
			        3393 => x"00000000",		-- colors: 40, 40, 40, 40
			        3394 => x"00000000",		-- colors: 40, 40, 40, 40
			        3395 => x"00000000",		-- colors: 40, 40, 40, 40
			        3396 => x"00000000",		-- colors: 40, 40, 40, 40
			        3397 => x"00000000",		-- colors: 40, 40, 40, 40
			        3398 => x"00000000",		-- colors: 40, 40, 40, 40
			        3399 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3400 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3401 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3402 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3403 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3404 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3405 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3406 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3407 => x"00000000",		-- colors: 40, 40, 40, 40
			        3408 => x"00000000",		-- colors: 40, 40, 40, 40
			        3409 => x"00000000",		-- colors: 40, 40, 40, 40
			        3410 => x"00000000",		-- colors: 40, 40, 40, 40
			        3411 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3412 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3413 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3414 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3415 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3416 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3417 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3418 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3419 => x"00000000",		-- colors: 40, 40, 40, 40
			        3420 => x"00000000",		-- colors: 40, 40, 40, 40
			        3421 => x"00000000",		-- colors: 40, 40, 40, 40
			        3422 => x"00000000",		-- colors: 40, 40, 40, 40
			        3423 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3424 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3425 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3426 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3427 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3428 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3429 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3430 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3431 => x"00000000",		-- colors: 40, 40, 40, 40
			        3432 => x"00000000",		-- colors: 40, 40, 40, 40
			        3433 => x"00000000",		-- colors: 40, 40, 40, 40
			        3434 => x"00000000",		-- colors: 40, 40, 40, 40
			        3435 => x"00000000",		-- colors: 40, 40, 40, 40
			        3436 => x"00000000",		-- colors: 40, 40, 40, 40
			        3437 => x"00000000",		-- colors: 40, 40, 40, 40
			        3438 => x"00000000",		-- colors: 40, 40, 40, 40
			        3439 => x"00000000",		-- colors: 40, 40, 40, 40
			        3440 => x"00000000",		-- colors: 40, 40, 40, 40
			        3441 => x"00000000",		-- colors: 40, 40, 40, 40
			        3442 => x"00000000",		-- colors: 40, 40, 40, 40
			        3443 => x"00000000",		-- colors: 40, 40, 40, 40
			        3444 => x"00000000",		-- colors: 40, 40, 40, 40
			        3445 => x"00000000",		-- colors: 40, 40, 40, 40
			        3446 => x"00000000",		-- colors: 40, 40, 40, 40
			        3447 => x"00000000",		-- colors: 40, 40, 40, 40
			        3448 => x"00000000",		-- colors: 40, 40, 40, 40
			        3449 => x"00000000",		-- colors: 40, 40, 40, 40
			        3450 => x"00000000",		-- colors: 40, 40, 40, 40
			        3451 => x"00000000",		-- colors: 40, 40, 40, 40
			        3452 => x"00000000",		-- colors: 40, 40, 40, 40
			        3453 => x"00000000",		-- colors: 40, 40, 40, 40
			        3454 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 50
			        3455 => x"00000000",		-- colors: 40, 40, 40, 40
			        3456 => x"00000000",		-- colors: 40, 40, 40, 40
			        3457 => x"00000000",		-- colors: 40, 40, 40, 40
			        3458 => x"00000000",		-- colors: 40, 40, 40, 40
			        3459 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3460 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3461 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3462 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3463 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3464 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3465 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3466 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3467 => x"00000000",		-- colors: 40, 40, 40, 40
			        3468 => x"00000000",		-- colors: 40, 40, 40, 40
			        3469 => x"00000000",		-- colors: 40, 40, 40, 40
			        3470 => x"00000000",		-- colors: 40, 40, 40, 40
			        3471 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3472 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3473 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3474 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3475 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3476 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3477 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3478 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3479 => x"00000000",		-- colors: 40, 40, 40, 40
			        3480 => x"00000000",		-- colors: 40, 40, 40, 40
			        3481 => x"00000000",		-- colors: 40, 40, 40, 40
			        3482 => x"00000000",		-- colors: 40, 40, 40, 40
			        3483 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3484 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3485 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3486 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3487 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3488 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3489 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3490 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3491 => x"00000000",		-- colors: 40, 40, 40, 40
			        3492 => x"00000000",		-- colors: 40, 40, 40, 40
			        3493 => x"00000000",		-- colors: 40, 40, 40, 40
			        3494 => x"00000000",		-- colors: 40, 40, 40, 40
			        3495 => x"32323232",		-- colors: 50, 50, 50, 50
			        3496 => x"32323232",		-- colors: 50, 50, 50, 50
			        3497 => x"32323232",		-- colors: 50, 50, 50, 50
			        3498 => x"32323232",		-- colors: 50, 50, 50, 50
			        3499 => x"00000000",		-- colors: 40, 40, 40, 40
			        3500 => x"00000000",		-- colors: 40, 40, 40, 40
			        3501 => x"00000000",		-- colors: 40, 40, 40, 40
			        3502 => x"00000000",		-- colors: 40, 40, 40, 40
			        3503 => x"00000000",		-- colors: 40, 40, 40, 40
			        3504 => x"00000000",		-- colors: 40, 40, 40, 40
			        3505 => x"00000000",		-- colors: 40, 40, 40, 40
			        3506 => x"00000000",		-- colors: 40, 40, 40, 40
			        3507 => x"00000000",		-- colors: 40, 40, 40, 40
			        3508 => x"00000000",		-- colors: 40, 40, 40, 40
			        3509 => x"00000000",		-- colors: 40, 40, 40, 40
			        3510 => x"00000000",		-- colors: 40, 40, 40, 40
			        3511 => x"32323232",		-- colors: 50, 50, 50, 50
			        3512 => x"32323232",		-- colors: 50, 50, 50, 50
			        3513 => x"32323232",		-- colors: 50, 50, 50, 50
			        3514 => x"32323232",		-- colors: 50, 50, 50, 50
			        3515 => x"00000000",		-- colors: 40, 40, 40, 40
			        3516 => x"00000000",		-- colors: 40, 40, 40, 40
			        3517 => x"00000000",		-- colors: 40, 40, 40, 40
			        3518 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 51
			        3519 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3520 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3521 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3522 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3523 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3524 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3525 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3526 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3527 => x"00000000",		-- colors: 40, 40, 40, 40
			        3528 => x"00000000",		-- colors: 40, 40, 40, 40
			        3529 => x"00000000",		-- colors: 40, 40, 40, 40
			        3530 => x"00000000",		-- colors: 40, 40, 40, 40
			        3531 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3532 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3533 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3534 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3535 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3536 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3537 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3538 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3539 => x"00000000",		-- colors: 40, 40, 40, 40
			        3540 => x"00000000",		-- colors: 40, 40, 40, 40
			        3541 => x"00000000",		-- colors: 40, 40, 40, 40
			        3542 => x"00000000",		-- colors: 40, 40, 40, 40
			        3543 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3544 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3545 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3546 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3547 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3548 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3549 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3550 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3551 => x"00000000",		-- colors: 40, 40, 40, 40
			        3552 => x"00000000",		-- colors: 40, 40, 40, 40
			        3553 => x"00000000",		-- colors: 40, 40, 40, 40
			        3554 => x"00000000",		-- colors: 40, 40, 40, 40
			        3555 => x"00000000",		-- colors: 40, 40, 40, 40
			        3556 => x"00000000",		-- colors: 40, 40, 40, 40
			        3557 => x"00000000",		-- colors: 40, 40, 40, 40
			        3558 => x"00000000",		-- colors: 40, 40, 40, 40
			        3559 => x"00000000",		-- colors: 40, 40, 40, 40
			        3560 => x"00000000",		-- colors: 40, 40, 40, 40
			        3561 => x"00000000",		-- colors: 40, 40, 40, 40
			        3562 => x"00000000",		-- colors: 40, 40, 40, 40
			        3563 => x"00000000",		-- colors: 40, 40, 40, 40
			        3564 => x"00000000",		-- colors: 40, 40, 40, 40
			        3565 => x"00000000",		-- colors: 40, 40, 40, 40
			        3566 => x"00000000",		-- colors: 40, 40, 40, 40
			        3567 => x"00000000",		-- colors: 40, 40, 40, 40
			        3568 => x"00000000",		-- colors: 40, 40, 40, 40
			        3569 => x"00000000",		-- colors: 40, 40, 40, 40
			        3570 => x"00000000",		-- colors: 40, 40, 40, 40
			        3571 => x"00000000",		-- colors: 40, 40, 40, 40
			        3572 => x"00000000",		-- colors: 40, 40, 40, 40
			        3573 => x"00000000",		-- colors: 40, 40, 40, 40
			        3574 => x"00000000",		-- colors: 40, 40, 40, 40
			        3575 => x"00000000",		-- colors: 40, 40, 40, 40
			        3576 => x"00000000",		-- colors: 40, 40, 40, 40
			        3577 => x"00000000",		-- colors: 40, 40, 40, 40
			        3578 => x"00000000",		-- colors: 40, 40, 40, 40
			        3579 => x"00000000",		-- colors: 40, 40, 40, 40
			        3580 => x"00000000",		-- colors: 40, 40, 40, 40
			        3581 => x"00000000",		-- colors: 40, 40, 40, 40
			        3582 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 52
			        3583 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3584 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3585 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3586 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3587 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3588 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3589 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3590 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3591 => x"00000000",		-- colors: 40, 40, 40, 40
			        3592 => x"00000000",		-- colors: 40, 40, 40, 40
			        3593 => x"00000000",		-- colors: 40, 40, 40, 40
			        3594 => x"00000000",		-- colors: 40, 40, 40, 40
			        3595 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3596 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3597 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3598 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3599 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3600 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3601 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3602 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3603 => x"00000000",		-- colors: 40, 40, 40, 40
			        3604 => x"00000000",		-- colors: 40, 40, 40, 40
			        3605 => x"00000000",		-- colors: 40, 40, 40, 40
			        3606 => x"00000000",		-- colors: 40, 40, 40, 40
			        3607 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3608 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3609 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3610 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3611 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3612 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3613 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3614 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3615 => x"00000000",		-- colors: 40, 40, 40, 40
			        3616 => x"00000000",		-- colors: 40, 40, 40, 40
			        3617 => x"00000000",		-- colors: 40, 40, 40, 40
			        3618 => x"00000000",		-- colors: 40, 40, 40, 40
			        3619 => x"00000000",		-- colors: 40, 40, 40, 40
			        3620 => x"00000000",		-- colors: 40, 40, 40, 40
			        3621 => x"00000000",		-- colors: 40, 40, 40, 40
			        3622 => x"00000000",		-- colors: 40, 40, 40, 40
			        3623 => x"00000000",		-- colors: 40, 40, 40, 40
			        3624 => x"00000000",		-- colors: 40, 40, 40, 40
			        3625 => x"00000000",		-- colors: 40, 40, 40, 40
			        3626 => x"00000000",		-- colors: 40, 40, 40, 40
			        3627 => x"00000000",		-- colors: 40, 40, 40, 40
			        3628 => x"00000000",		-- colors: 40, 40, 40, 40
			        3629 => x"00000000",		-- colors: 40, 40, 40, 40
			        3630 => x"00000000",		-- colors: 40, 40, 40, 40
			        3631 => x"00000000",		-- colors: 40, 40, 40, 40
			        3632 => x"00000000",		-- colors: 40, 40, 40, 40
			        3633 => x"00000000",		-- colors: 40, 40, 40, 40
			        3634 => x"00000000",		-- colors: 40, 40, 40, 40
			        3635 => x"00000000",		-- colors: 40, 40, 40, 40
			        3636 => x"00000000",		-- colors: 40, 40, 40, 40
			        3637 => x"00000000",		-- colors: 40, 40, 40, 40
			        3638 => x"00000000",		-- colors: 40, 40, 40, 40
			        3639 => x"00000000",		-- colors: 40, 40, 40, 40
			        3640 => x"00000000",		-- colors: 40, 40, 40, 40
			        3641 => x"00000000",		-- colors: 40, 40, 40, 40
			        3642 => x"00000000",		-- colors: 40, 40, 40, 40
			        3643 => x"00000000",		-- colors: 40, 40, 40, 40
			        3644 => x"00000000",		-- colors: 40, 40, 40, 40
			        3645 => x"00000000",		-- colors: 40, 40, 40, 40
			        3646 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 53
			        3647 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3648 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3649 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3650 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3651 => x"00000000",		-- colors: 40, 40, 40, 40
			        3652 => x"00000000",		-- colors: 40, 40, 40, 40
			        3653 => x"00000000",		-- colors: 40, 40, 40, 40
			        3654 => x"00000000",		-- colors: 40, 40, 40, 40
			        3655 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3656 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3657 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3658 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3659 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3660 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3661 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3662 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3663 => x"00000000",		-- colors: 40, 40, 40, 40
			        3664 => x"00000000",		-- colors: 40, 40, 40, 40
			        3665 => x"00000000",		-- colors: 40, 40, 40, 40
			        3666 => x"00000000",		-- colors: 40, 40, 40, 40
			        3667 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3668 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3669 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3670 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3671 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3672 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3673 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3674 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3675 => x"00000000",		-- colors: 40, 40, 40, 40
			        3676 => x"00000000",		-- colors: 40, 40, 40, 40
			        3677 => x"00000000",		-- colors: 40, 40, 40, 40
			        3678 => x"00000000",		-- colors: 40, 40, 40, 40
			        3679 => x"00000000",		-- colors: 40, 40, 40, 40
			        3680 => x"00000000",		-- colors: 40, 40, 40, 40
			        3681 => x"00000000",		-- colors: 40, 40, 40, 40
			        3682 => x"00000000",		-- colors: 40, 40, 40, 40
			        3683 => x"00000000",		-- colors: 40, 40, 40, 40
			        3684 => x"00000000",		-- colors: 40, 40, 40, 40
			        3685 => x"00000000",		-- colors: 40, 40, 40, 40
			        3686 => x"00000000",		-- colors: 40, 40, 40, 40
			        3687 => x"00000000",		-- colors: 40, 40, 40, 40
			        3688 => x"00000000",		-- colors: 40, 40, 40, 40
			        3689 => x"00000000",		-- colors: 40, 40, 40, 40
			        3690 => x"00000000",		-- colors: 40, 40, 40, 40
			        3691 => x"00000000",		-- colors: 40, 40, 40, 40
			        3692 => x"00000000",		-- colors: 40, 40, 40, 40
			        3693 => x"00000000",		-- colors: 40, 40, 40, 40
			        3694 => x"00000000",		-- colors: 40, 40, 40, 40
			        3695 => x"00000000",		-- colors: 40, 40, 40, 40
			        3696 => x"00000000",		-- colors: 40, 40, 40, 40
			        3697 => x"00000000",		-- colors: 40, 40, 40, 40
			        3698 => x"00000000",		-- colors: 40, 40, 40, 40
			        3699 => x"00000000",		-- colors: 40, 40, 40, 40
			        3700 => x"00000000",		-- colors: 40, 40, 40, 40
			        3701 => x"00000000",		-- colors: 40, 40, 40, 40
			        3702 => x"00000000",		-- colors: 40, 40, 40, 40
			        3703 => x"00000000",		-- colors: 40, 40, 40, 40
			        3704 => x"00000000",		-- colors: 40, 40, 40, 40
			        3705 => x"00000000",		-- colors: 40, 40, 40, 40
			        3706 => x"00000000",		-- colors: 40, 40, 40, 40
			        3707 => x"00000000",		-- colors: 40, 40, 40, 40
			        3708 => x"00000000",		-- colors: 40, 40, 40, 40
			        3709 => x"00000000",		-- colors: 40, 40, 40, 40
			        3710 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 54
			        3711 => x"00000000",		-- colors: 40, 40, 40, 40
			        3712 => x"00000000",		-- colors: 40, 40, 40, 40
			        3713 => x"00000000",		-- colors: 40, 40, 40, 40
			        3714 => x"00000000",		-- colors: 40, 40, 40, 40
			        3715 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3716 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3717 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3718 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3719 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3720 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3721 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3722 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3723 => x"00000000",		-- colors: 40, 40, 40, 40
			        3724 => x"00000000",		-- colors: 40, 40, 40, 40
			        3725 => x"00000000",		-- colors: 40, 40, 40, 40
			        3726 => x"00000000",		-- colors: 40, 40, 40, 40
			        3727 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3728 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3729 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3730 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3731 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3732 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3733 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3734 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3735 => x"00000000",		-- colors: 40, 40, 40, 40
			        3736 => x"00000000",		-- colors: 40, 40, 40, 40
			        3737 => x"00000000",		-- colors: 40, 40, 40, 40
			        3738 => x"00000000",		-- colors: 40, 40, 40, 40
			        3739 => x"00000000",		-- colors: 40, 40, 40, 40
			        3740 => x"00000000",		-- colors: 40, 40, 40, 40
			        3741 => x"00000000",		-- colors: 40, 40, 40, 40
			        3742 => x"00000000",		-- colors: 40, 40, 40, 40
			        3743 => x"00000000",		-- colors: 40, 40, 40, 40
			        3744 => x"00000000",		-- colors: 40, 40, 40, 40
			        3745 => x"00000000",		-- colors: 40, 40, 40, 40
			        3746 => x"00000000",		-- colors: 40, 40, 40, 40
			        3747 => x"00000000",		-- colors: 40, 40, 40, 40
			        3748 => x"00000000",		-- colors: 40, 40, 40, 40
			        3749 => x"00000000",		-- colors: 40, 40, 40, 40
			        3750 => x"00000000",		-- colors: 40, 40, 40, 40
			        3751 => x"00000000",		-- colors: 40, 40, 40, 40
			        3752 => x"00000000",		-- colors: 40, 40, 40, 40
			        3753 => x"00000000",		-- colors: 40, 40, 40, 40
			        3754 => x"00000000",		-- colors: 40, 40, 40, 40
			        3755 => x"00000000",		-- colors: 40, 40, 40, 40
			        3756 => x"00000000",		-- colors: 40, 40, 40, 40
			        3757 => x"00000000",		-- colors: 40, 40, 40, 40
			        3758 => x"00000000",		-- colors: 40, 40, 40, 40
			        3759 => x"00000000",		-- colors: 40, 40, 40, 40
			        3760 => x"00000000",		-- colors: 40, 40, 40, 40
			        3761 => x"00000000",		-- colors: 40, 40, 40, 40
			        3762 => x"00000000",		-- colors: 40, 40, 40, 40
			        3763 => x"00000000",		-- colors: 40, 40, 40, 40
			        3764 => x"00000000",		-- colors: 40, 40, 40, 40
			        3765 => x"00000000",		-- colors: 40, 40, 40, 40
			        3766 => x"00000000",		-- colors: 40, 40, 40, 40
			        3767 => x"00000000",		-- colors: 40, 40, 40, 40
			        3768 => x"00000000",		-- colors: 40, 40, 40, 40
			        3769 => x"00000000",		-- colors: 40, 40, 40, 40
			        3770 => x"00000000",		-- colors: 40, 40, 40, 40
			        3771 => x"00000000",		-- colors: 40, 40, 40, 40
			        3772 => x"00000000",		-- colors: 40, 40, 40, 40
			        3773 => x"00000000",		-- colors: 40, 40, 40, 40
			        3774 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 55
			        3775 => x"00000000",		-- colors: 40, 40, 40, 40
			        3776 => x"00000000",		-- colors: 40, 40, 40, 40
			        3777 => x"00000000",		-- colors: 40, 40, 40, 40
			        3778 => x"00000000",		-- colors: 40, 40, 40, 40
			        3779 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3780 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3781 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3782 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3783 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3784 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3785 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3786 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3787 => x"00000000",		-- colors: 40, 40, 40, 40
			        3788 => x"00000000",		-- colors: 40, 40, 40, 40
			        3789 => x"00000000",		-- colors: 40, 40, 40, 40
			        3790 => x"00000000",		-- colors: 40, 40, 40, 40
			        3791 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3792 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3793 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3794 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3795 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3796 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3797 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3798 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3799 => x"00000000",		-- colors: 40, 40, 40, 40
			        3800 => x"00000000",		-- colors: 40, 40, 40, 40
			        3801 => x"00000000",		-- colors: 40, 40, 40, 40
			        3802 => x"00000000",		-- colors: 40, 40, 40, 40
			        3803 => x"00000000",		-- colors: 40, 40, 40, 40
			        3804 => x"00000000",		-- colors: 40, 40, 40, 40
			        3805 => x"00000000",		-- colors: 40, 40, 40, 40
			        3806 => x"00000000",		-- colors: 40, 40, 40, 40
			        3807 => x"00000000",		-- colors: 40, 40, 40, 40
			        3808 => x"00000000",		-- colors: 40, 40, 40, 40
			        3809 => x"00000000",		-- colors: 40, 40, 40, 40
			        3810 => x"00000000",		-- colors: 40, 40, 40, 40
			        3811 => x"00000000",		-- colors: 40, 40, 40, 40
			        3812 => x"00000000",		-- colors: 40, 40, 40, 40
			        3813 => x"00000000",		-- colors: 40, 40, 40, 40
			        3814 => x"00000000",		-- colors: 40, 40, 40, 40
			        3815 => x"00000000",		-- colors: 40, 40, 40, 40
			        3816 => x"00000000",		-- colors: 40, 40, 40, 40
			        3817 => x"00000000",		-- colors: 40, 40, 40, 40
			        3818 => x"00000000",		-- colors: 40, 40, 40, 40
			        3819 => x"00000000",		-- colors: 40, 40, 40, 40
			        3820 => x"00000000",		-- colors: 40, 40, 40, 40
			        3821 => x"00000000",		-- colors: 40, 40, 40, 40
			        3822 => x"00000000",		-- colors: 40, 40, 40, 40
			        3823 => x"00000000",		-- colors: 40, 40, 40, 40
			        3824 => x"00000000",		-- colors: 40, 40, 40, 40
			        3825 => x"00000000",		-- colors: 40, 40, 40, 40
			        3826 => x"00000000",		-- colors: 40, 40, 40, 40
			        3827 => x"00000000",		-- colors: 40, 40, 40, 40
			        3828 => x"00000000",		-- colors: 40, 40, 40, 40
			        3829 => x"00000000",		-- colors: 40, 40, 40, 40
			        3830 => x"00000000",		-- colors: 40, 40, 40, 40
			        3831 => x"00000000",		-- colors: 40, 40, 40, 40
			        3832 => x"00000000",		-- colors: 40, 40, 40, 40
			        3833 => x"00000000",		-- colors: 40, 40, 40, 40
			        3834 => x"00000000",		-- colors: 40, 40, 40, 40
			        3835 => x"00000000",		-- colors: 40, 40, 40, 40
			        3836 => x"00000000",		-- colors: 40, 40, 40, 40
			        3837 => x"00000000",		-- colors: 40, 40, 40, 40
			        3838 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 56
			        3839 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3840 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3841 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3842 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3843 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3844 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3845 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3846 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3847 => x"00000000",		-- colors: 40, 40, 40, 40
			        3848 => x"00000000",		-- colors: 40, 40, 40, 40
			        3849 => x"00000000",		-- colors: 40, 40, 40, 40
			        3850 => x"00000000",		-- colors: 40, 40, 40, 40
			        3851 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3852 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3853 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3854 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3855 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3856 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3857 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3858 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3859 => x"00000000",		-- colors: 40, 40, 40, 40
			        3860 => x"00000000",		-- colors: 40, 40, 40, 40
			        3861 => x"00000000",		-- colors: 40, 40, 40, 40
			        3862 => x"00000000",		-- colors: 40, 40, 40, 40
			        3863 => x"32323232",		-- colors: 50, 50, 50, 50
			        3864 => x"32323232",		-- colors: 50, 50, 50, 50
			        3865 => x"32323232",		-- colors: 50, 50, 50, 50
			        3866 => x"32323232",		-- colors: 50, 50, 50, 50
			        3867 => x"00000000",		-- colors: 40, 40, 40, 40
			        3868 => x"00000000",		-- colors: 40, 40, 40, 40
			        3869 => x"00000000",		-- colors: 40, 40, 40, 40
			        3870 => x"00000000",		-- colors: 40, 40, 40, 40
			        3871 => x"00000000",		-- colors: 40, 40, 40, 40
			        3872 => x"00000000",		-- colors: 40, 40, 40, 40
			        3873 => x"00000000",		-- colors: 40, 40, 40, 40
			        3874 => x"00000000",		-- colors: 40, 40, 40, 40
			        3875 => x"00000000",		-- colors: 40, 40, 40, 40
			        3876 => x"00000000",		-- colors: 40, 40, 40, 40
			        3877 => x"00000000",		-- colors: 40, 40, 40, 40
			        3878 => x"00000000",		-- colors: 40, 40, 40, 40
			        3879 => x"00000000",		-- colors: 40, 40, 40, 40
			        3880 => x"00000000",		-- colors: 40, 40, 40, 40
			        3881 => x"00000000",		-- colors: 40, 40, 40, 40
			        3882 => x"00000000",		-- colors: 40, 40, 40, 40
			        3883 => x"00000000",		-- colors: 40, 40, 40, 40
			        3884 => x"00000000",		-- colors: 40, 40, 40, 40
			        3885 => x"00000000",		-- colors: 40, 40, 40, 40
			        3886 => x"00000000",		-- colors: 40, 40, 40, 40
			        3887 => x"00000000",		-- colors: 40, 40, 40, 40
			        3888 => x"00000000",		-- colors: 40, 40, 40, 40
			        3889 => x"00000000",		-- colors: 40, 40, 40, 40
			        3890 => x"00000000",		-- colors: 40, 40, 40, 40
			        3891 => x"00000000",		-- colors: 40, 40, 40, 40
			        3892 => x"00000000",		-- colors: 40, 40, 40, 40
			        3893 => x"00000000",		-- colors: 40, 40, 40, 40
			        3894 => x"00000000",		-- colors: 40, 40, 40, 40
			        3895 => x"00000000",		-- colors: 40, 40, 40, 40
			        3896 => x"00000000",		-- colors: 40, 40, 40, 40
			        3897 => x"00000000",		-- colors: 40, 40, 40, 40
			        3898 => x"00000000",		-- colors: 40, 40, 40, 40
			        3899 => x"00000000",		-- colors: 40, 40, 40, 40
			        3900 => x"00000000",		-- colors: 40, 40, 40, 40
			        3901 => x"00000000",		-- colors: 40, 40, 40, 40
			        3902 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 57
			        3903 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3904 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3905 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3906 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3907 => x"00000000",		-- colors: 40, 40, 40, 40
			        3908 => x"00000000",		-- colors: 40, 40, 40, 40
			        3909 => x"00000000",		-- colors: 40, 40, 40, 40
			        3910 => x"00000000",		-- colors: 40, 40, 40, 40
			        3911 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3912 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3913 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3914 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3915 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3916 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3917 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3918 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3919 => x"00000000",		-- colors: 40, 40, 40, 40
			        3920 => x"00000000",		-- colors: 40, 40, 40, 40
			        3921 => x"00000000",		-- colors: 40, 40, 40, 40
			        3922 => x"00000000",		-- colors: 40, 40, 40, 40
			        3923 => x"00000000",		-- colors: 40, 40, 40, 40
			        3924 => x"00000000",		-- colors: 40, 40, 40, 40
			        3925 => x"00000000",		-- colors: 40, 40, 40, 40
			        3926 => x"00000000",		-- colors: 40, 40, 40, 40
			        3927 => x"00000000",		-- colors: 40, 40, 40, 40
			        3928 => x"00000000",		-- colors: 40, 40, 40, 40
			        3929 => x"00000000",		-- colors: 40, 40, 40, 40
			        3930 => x"00000000",		-- colors: 40, 40, 40, 40
			        3931 => x"00000000",		-- colors: 40, 40, 40, 40
			        3932 => x"00000000",		-- colors: 40, 40, 40, 40
			        3933 => x"00000000",		-- colors: 40, 40, 40, 40
			        3934 => x"00000000",		-- colors: 40, 40, 40, 40
			        3935 => x"00000000",		-- colors: 40, 40, 40, 40
			        3936 => x"00000000",		-- colors: 40, 40, 40, 40
			        3937 => x"00000000",		-- colors: 40, 40, 40, 40
			        3938 => x"00000000",		-- colors: 40, 40, 40, 40
			        3939 => x"00000000",		-- colors: 40, 40, 40, 40
			        3940 => x"00000000",		-- colors: 40, 40, 40, 40
			        3941 => x"00000000",		-- colors: 40, 40, 40, 40
			        3942 => x"00000000",		-- colors: 40, 40, 40, 40
			        3943 => x"00000000",		-- colors: 40, 40, 40, 40
			        3944 => x"00000000",		-- colors: 40, 40, 40, 40
			        3945 => x"00000000",		-- colors: 40, 40, 40, 40
			        3946 => x"00000000",		-- colors: 40, 40, 40, 40
			        3947 => x"00000000",		-- colors: 40, 40, 40, 40
			        3948 => x"00000000",		-- colors: 40, 40, 40, 40
			        3949 => x"00000000",		-- colors: 40, 40, 40, 40
			        3950 => x"00000000",		-- colors: 40, 40, 40, 40
			        3951 => x"00000000",		-- colors: 40, 40, 40, 40
			        3952 => x"00000000",		-- colors: 40, 40, 40, 40
			        3953 => x"00000000",		-- colors: 40, 40, 40, 40
			        3954 => x"00000000",		-- colors: 40, 40, 40, 40
			        3955 => x"00000000",		-- colors: 40, 40, 40, 40
			        3956 => x"00000000",		-- colors: 40, 40, 40, 40
			        3957 => x"00000000",		-- colors: 40, 40, 40, 40
			        3958 => x"00000000",		-- colors: 40, 40, 40, 40
			        3959 => x"00000000",		-- colors: 40, 40, 40, 40
			        3960 => x"00000000",		-- colors: 40, 40, 40, 40
			        3961 => x"00000000",		-- colors: 40, 40, 40, 40
			        3962 => x"00000000",		-- colors: 40, 40, 40, 40
			        3963 => x"00000000",		-- colors: 40, 40, 40, 40
			        3964 => x"00000000",		-- colors: 40, 40, 40, 40
			        3965 => x"00000000",		-- colors: 40, 40, 40, 40
			        3966 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 58
			        3967 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3968 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3969 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3970 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3971 => x"00000000",		-- colors: 40, 40, 40, 40
			        3972 => x"00000000",		-- colors: 40, 40, 40, 40
			        3973 => x"00000000",		-- colors: 40, 40, 40, 40
			        3974 => x"00000000",		-- colors: 40, 40, 40, 40
			        3975 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3976 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3977 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3978 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3979 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3980 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3981 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3982 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        3983 => x"00000000",		-- colors: 40, 40, 40, 40
			        3984 => x"00000000",		-- colors: 40, 40, 40, 40
			        3985 => x"00000000",		-- colors: 40, 40, 40, 40
			        3986 => x"00000000",		-- colors: 40, 40, 40, 40
			        3987 => x"00000000",		-- colors: 40, 40, 40, 40
			        3988 => x"00000000",		-- colors: 40, 40, 40, 40
			        3989 => x"00000000",		-- colors: 40, 40, 40, 40
			        3990 => x"00000000",		-- colors: 40, 40, 40, 40
			        3991 => x"00000000",		-- colors: 40, 40, 40, 40
			        3992 => x"00000000",		-- colors: 40, 40, 40, 40
			        3993 => x"00000000",		-- colors: 40, 40, 40, 40
			        3994 => x"00000000",		-- colors: 40, 40, 40, 40
			        3995 => x"00000000",		-- colors: 40, 40, 40, 40
			        3996 => x"00000000",		-- colors: 40, 40, 40, 40
			        3997 => x"00000000",		-- colors: 40, 40, 40, 40
			        3998 => x"00000000",		-- colors: 40, 40, 40, 40
			        3999 => x"00000000",		-- colors: 40, 40, 40, 40
			        4000 => x"00000000",		-- colors: 40, 40, 40, 40
			        4001 => x"00000000",		-- colors: 40, 40, 40, 40
			        4002 => x"00000000",		-- colors: 40, 40, 40, 40
			        4003 => x"00000000",		-- colors: 40, 40, 40, 40
			        4004 => x"00000000",		-- colors: 40, 40, 40, 40
			        4005 => x"00000000",		-- colors: 40, 40, 40, 40
			        4006 => x"00000000",		-- colors: 40, 40, 40, 40
			        4007 => x"00000000",		-- colors: 40, 40, 40, 40
			        4008 => x"00000000",		-- colors: 40, 40, 40, 40
			        4009 => x"00000000",		-- colors: 40, 40, 40, 40
			        4010 => x"00000000",		-- colors: 40, 40, 40, 40
			        4011 => x"00000000",		-- colors: 40, 40, 40, 40
			        4012 => x"00000000",		-- colors: 40, 40, 40, 40
			        4013 => x"00000000",		-- colors: 40, 40, 40, 40
			        4014 => x"00000000",		-- colors: 40, 40, 40, 40
			        4015 => x"00000000",		-- colors: 40, 40, 40, 40
			        4016 => x"00000000",		-- colors: 40, 40, 40, 40
			        4017 => x"00000000",		-- colors: 40, 40, 40, 40
			        4018 => x"00000000",		-- colors: 40, 40, 40, 40
			        4019 => x"00000000",		-- colors: 40, 40, 40, 40
			        4020 => x"00000000",		-- colors: 40, 40, 40, 40
			        4021 => x"00000000",		-- colors: 40, 40, 40, 40
			        4022 => x"00000000",		-- colors: 40, 40, 40, 40
			        4023 => x"00000000",		-- colors: 40, 40, 40, 40
			        4024 => x"00000000",		-- colors: 40, 40, 40, 40
			        4025 => x"00000000",		-- colors: 40, 40, 40, 40
			        4026 => x"00000000",		-- colors: 40, 40, 40, 40
			        4027 => x"00000000",		-- colors: 40, 40, 40, 40
			        4028 => x"00000000",		-- colors: 40, 40, 40, 40
			        4029 => x"00000000",		-- colors: 40, 40, 40, 40
			        4030 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 59
			        4031 => x"00000000",		-- colors: 40, 40, 40, 40
			        4032 => x"00000000",		-- colors: 40, 40, 40, 40
			        4033 => x"00000000",		-- colors: 40, 40, 40, 40
			        4034 => x"00000000",		-- colors: 40, 40, 40, 40
			        4035 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4036 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4037 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4038 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4039 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4040 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4041 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4042 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4043 => x"00000000",		-- colors: 40, 40, 40, 40
			        4044 => x"00000000",		-- colors: 40, 40, 40, 40
			        4045 => x"00000000",		-- colors: 40, 40, 40, 40
			        4046 => x"00000000",		-- colors: 40, 40, 40, 40
			        4047 => x"00000000",		-- colors: 40, 40, 40, 40
			        4048 => x"00000000",		-- colors: 40, 40, 40, 40
			        4049 => x"00000000",		-- colors: 40, 40, 40, 40
			        4050 => x"00000000",		-- colors: 40, 40, 40, 40
			        4051 => x"00000000",		-- colors: 40, 40, 40, 40
			        4052 => x"00000000",		-- colors: 40, 40, 40, 40
			        4053 => x"00000000",		-- colors: 40, 40, 40, 40
			        4054 => x"00000000",		-- colors: 40, 40, 40, 40
			        4055 => x"00000000",		-- colors: 40, 40, 40, 40
			        4056 => x"00000000",		-- colors: 40, 40, 40, 40
			        4057 => x"00000000",		-- colors: 40, 40, 40, 40
			        4058 => x"00000000",		-- colors: 40, 40, 40, 40
			        4059 => x"00000000",		-- colors: 40, 40, 40, 40
			        4060 => x"00000000",		-- colors: 40, 40, 40, 40
			        4061 => x"00000000",		-- colors: 40, 40, 40, 40
			        4062 => x"00000000",		-- colors: 40, 40, 40, 40
			        4063 => x"00000000",		-- colors: 40, 40, 40, 40
			        4064 => x"00000000",		-- colors: 40, 40, 40, 40
			        4065 => x"00000000",		-- colors: 40, 40, 40, 40
			        4066 => x"00000000",		-- colors: 40, 40, 40, 40
			        4067 => x"00000000",		-- colors: 40, 40, 40, 40
			        4068 => x"00000000",		-- colors: 40, 40, 40, 40
			        4069 => x"00000000",		-- colors: 40, 40, 40, 40
			        4070 => x"00000000",		-- colors: 40, 40, 40, 40
			        4071 => x"00000000",		-- colors: 40, 40, 40, 40
			        4072 => x"00000000",		-- colors: 40, 40, 40, 40
			        4073 => x"00000000",		-- colors: 40, 40, 40, 40
			        4074 => x"00000000",		-- colors: 40, 40, 40, 40
			        4075 => x"00000000",		-- colors: 40, 40, 40, 40
			        4076 => x"00000000",		-- colors: 40, 40, 40, 40
			        4077 => x"00000000",		-- colors: 40, 40, 40, 40
			        4078 => x"00000000",		-- colors: 40, 40, 40, 40
			        4079 => x"00000000",		-- colors: 40, 40, 40, 40
			        4080 => x"00000000",		-- colors: 40, 40, 40, 40
			        4081 => x"00000000",		-- colors: 40, 40, 40, 40
			        4082 => x"00000000",		-- colors: 40, 40, 40, 40
			        4083 => x"00000000",		-- colors: 40, 40, 40, 40
			        4084 => x"00000000",		-- colors: 40, 40, 40, 40
			        4085 => x"00000000",		-- colors: 40, 40, 40, 40
			        4086 => x"00000000",		-- colors: 40, 40, 40, 40
			        4087 => x"00000000",		-- colors: 40, 40, 40, 40
			        4088 => x"00000000",		-- colors: 40, 40, 40, 40
			        4089 => x"00000000",		-- colors: 40, 40, 40, 40
			        4090 => x"00000000",		-- colors: 40, 40, 40, 40
			        4091 => x"00000000",		-- colors: 40, 40, 40, 40
			        4092 => x"00000000",		-- colors: 40, 40, 40, 40
			        4093 => x"00000000",		-- colors: 40, 40, 40, 40
			        4094 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 60
			        4095 => x"00000000",		-- colors: 40, 40, 40, 40
			        4096 => x"00000000",		-- colors: 40, 40, 40, 40
			        4097 => x"00000000",		-- colors: 40, 40, 40, 40
			        4098 => x"00000000",		-- colors: 40, 40, 40, 40
			        4099 => x"00000000",		-- colors: 40, 40, 40, 40
			        4100 => x"00000000",		-- colors: 40, 40, 40, 40
			        4101 => x"00000000",		-- colors: 40, 40, 40, 40
			        4102 => x"00000000",		-- colors: 40, 40, 40, 40
			        4103 => x"00000000",		-- colors: 40, 40, 40, 40
			        4104 => x"00000000",		-- colors: 40, 40, 40, 40
			        4105 => x"00000000",		-- colors: 40, 40, 40, 40
			        4106 => x"00000000",		-- colors: 40, 40, 40, 40
			        4107 => x"00000000",		-- colors: 40, 40, 40, 40
			        4108 => x"00000000",		-- colors: 40, 40, 40, 40
			        4109 => x"00000000",		-- colors: 40, 40, 40, 40
			        4110 => x"00000000",		-- colors: 40, 40, 40, 40
			        4111 => x"00000000",		-- colors: 40, 40, 40, 40
			        4112 => x"00000000",		-- colors: 40, 40, 40, 40
			        4113 => x"00000000",		-- colors: 40, 40, 40, 40
			        4114 => x"00000000",		-- colors: 40, 40, 40, 40
			        4115 => x"00000000",		-- colors: 40, 40, 40, 40
			        4116 => x"00000000",		-- colors: 40, 40, 40, 40
			        4117 => x"00000000",		-- colors: 40, 40, 40, 40
			        4118 => x"00000000",		-- colors: 40, 40, 40, 40
			        4119 => x"00000000",		-- colors: 40, 40, 40, 40
			        4120 => x"00000000",		-- colors: 40, 40, 40, 40
			        4121 => x"00000000",		-- colors: 40, 40, 40, 40
			        4122 => x"00000000",		-- colors: 40, 40, 40, 40
			        4123 => x"00000000",		-- colors: 40, 40, 40, 40
			        4124 => x"00000000",		-- colors: 40, 40, 40, 40
			        4125 => x"00000000",		-- colors: 40, 40, 40, 40
			        4126 => x"00000000",		-- colors: 40, 40, 40, 40
			        4127 => x"00000000",		-- colors: 40, 40, 40, 40
			        4128 => x"00000000",		-- colors: 40, 40, 40, 40
			        4129 => x"00000000",		-- colors: 40, 40, 40, 40
			        4130 => x"00000000",		-- colors: 40, 40, 40, 40
			        4131 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4132 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4133 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4134 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4135 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4136 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4137 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4138 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4139 => x"00000000",		-- colors: 40, 40, 40, 40
			        4140 => x"00000000",		-- colors: 40, 40, 40, 40
			        4141 => x"00000000",		-- colors: 40, 40, 40, 40
			        4142 => x"00000000",		-- colors: 40, 40, 40, 40
			        4143 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4144 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4145 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4146 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4147 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4148 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4149 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4150 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4151 => x"00000000",		-- colors: 40, 40, 40, 40
			        4152 => x"00000000",		-- colors: 40, 40, 40, 40
			        4153 => x"00000000",		-- colors: 40, 40, 40, 40
			        4154 => x"00000000",		-- colors: 40, 40, 40, 40
			        4155 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4156 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4157 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4158 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60

			                --  sprite 61
			        4159 => x"00000000",		-- colors: 40, 40, 40, 40
			        4160 => x"00000000",		-- colors: 40, 40, 40, 40
			        4161 => x"00000000",		-- colors: 40, 40, 40, 40
			        4162 => x"00000000",		-- colors: 40, 40, 40, 40
			        4163 => x"00000000",		-- colors: 40, 40, 40, 40
			        4164 => x"00000000",		-- colors: 40, 40, 40, 40
			        4165 => x"00000000",		-- colors: 40, 40, 40, 40
			        4166 => x"00000000",		-- colors: 40, 40, 40, 40
			        4167 => x"00000000",		-- colors: 40, 40, 40, 40
			        4168 => x"00000000",		-- colors: 40, 40, 40, 40
			        4169 => x"00000000",		-- colors: 40, 40, 40, 40
			        4170 => x"00000000",		-- colors: 40, 40, 40, 40
			        4171 => x"00000000",		-- colors: 40, 40, 40, 40
			        4172 => x"00000000",		-- colors: 40, 40, 40, 40
			        4173 => x"00000000",		-- colors: 40, 40, 40, 40
			        4174 => x"00000000",		-- colors: 40, 40, 40, 40
			        4175 => x"00000000",		-- colors: 40, 40, 40, 40
			        4176 => x"00000000",		-- colors: 40, 40, 40, 40
			        4177 => x"00000000",		-- colors: 40, 40, 40, 40
			        4178 => x"00000000",		-- colors: 40, 40, 40, 40
			        4179 => x"00000000",		-- colors: 40, 40, 40, 40
			        4180 => x"00000000",		-- colors: 40, 40, 40, 40
			        4181 => x"00000000",		-- colors: 40, 40, 40, 40
			        4182 => x"00000000",		-- colors: 40, 40, 40, 40
			        4183 => x"00000000",		-- colors: 40, 40, 40, 40
			        4184 => x"00000000",		-- colors: 40, 40, 40, 40
			        4185 => x"00000000",		-- colors: 40, 40, 40, 40
			        4186 => x"00000000",		-- colors: 40, 40, 40, 40
			        4187 => x"00000000",		-- colors: 40, 40, 40, 40
			        4188 => x"00000000",		-- colors: 40, 40, 40, 40
			        4189 => x"00000000",		-- colors: 40, 40, 40, 40
			        4190 => x"00000000",		-- colors: 40, 40, 40, 40
			        4191 => x"00000000",		-- colors: 40, 40, 40, 40
			        4192 => x"00000000",		-- colors: 40, 40, 40, 40
			        4193 => x"00000000",		-- colors: 40, 40, 40, 40
			        4194 => x"00000000",		-- colors: 40, 40, 40, 40
			        4195 => x"00000000",		-- colors: 40, 40, 40, 40
			        4196 => x"00000000",		-- colors: 40, 40, 40, 40
			        4197 => x"00000000",		-- colors: 40, 40, 40, 40
			        4198 => x"00000000",		-- colors: 40, 40, 40, 40
			        4199 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4200 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4201 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4202 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4203 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4204 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4205 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4206 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4207 => x"00000000",		-- colors: 40, 40, 40, 40
			        4208 => x"00000000",		-- colors: 40, 40, 40, 40
			        4209 => x"00000000",		-- colors: 40, 40, 40, 40
			        4210 => x"00000000",		-- colors: 40, 40, 40, 40
			        4211 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4212 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4213 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4214 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4215 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4216 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4217 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4218 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4219 => x"00000000",		-- colors: 40, 40, 40, 40
			        4220 => x"00000000",		-- colors: 40, 40, 40, 40
			        4221 => x"00000000",		-- colors: 40, 40, 40, 40
			        4222 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 62
			        4223 => x"00000000",		-- colors: 40, 40, 40, 40
			        4224 => x"00000000",		-- colors: 40, 40, 40, 40
			        4225 => x"00000000",		-- colors: 40, 40, 40, 40
			        4226 => x"00000000",		-- colors: 40, 40, 40, 40
			        4227 => x"00000000",		-- colors: 40, 40, 40, 40
			        4228 => x"00000000",		-- colors: 40, 40, 40, 40
			        4229 => x"00000000",		-- colors: 40, 40, 40, 40
			        4230 => x"00000000",		-- colors: 40, 40, 40, 40
			        4231 => x"00000000",		-- colors: 40, 40, 40, 40
			        4232 => x"00000000",		-- colors: 40, 40, 40, 40
			        4233 => x"00000000",		-- colors: 40, 40, 40, 40
			        4234 => x"00000000",		-- colors: 40, 40, 40, 40
			        4235 => x"00000000",		-- colors: 40, 40, 40, 40
			        4236 => x"00000000",		-- colors: 40, 40, 40, 40
			        4237 => x"00000000",		-- colors: 40, 40, 40, 40
			        4238 => x"00000000",		-- colors: 40, 40, 40, 40
			        4239 => x"00000000",		-- colors: 40, 40, 40, 40
			        4240 => x"00000000",		-- colors: 40, 40, 40, 40
			        4241 => x"00000000",		-- colors: 40, 40, 40, 40
			        4242 => x"00000000",		-- colors: 40, 40, 40, 40
			        4243 => x"00000000",		-- colors: 40, 40, 40, 40
			        4244 => x"00000000",		-- colors: 40, 40, 40, 40
			        4245 => x"00000000",		-- colors: 40, 40, 40, 40
			        4246 => x"00000000",		-- colors: 40, 40, 40, 40
			        4247 => x"00000000",		-- colors: 40, 40, 40, 40
			        4248 => x"00000000",		-- colors: 40, 40, 40, 40
			        4249 => x"00000000",		-- colors: 40, 40, 40, 40
			        4250 => x"00000000",		-- colors: 40, 40, 40, 40
			        4251 => x"00000000",		-- colors: 40, 40, 40, 40
			        4252 => x"00000000",		-- colors: 40, 40, 40, 40
			        4253 => x"00000000",		-- colors: 40, 40, 40, 40
			        4254 => x"00000000",		-- colors: 40, 40, 40, 40
			        4255 => x"00000000",		-- colors: 40, 40, 40, 40
			        4256 => x"00000000",		-- colors: 40, 40, 40, 40
			        4257 => x"00000000",		-- colors: 40, 40, 40, 40
			        4258 => x"00000000",		-- colors: 40, 40, 40, 40
			        4259 => x"00000000",		-- colors: 40, 40, 40, 40
			        4260 => x"00000000",		-- colors: 40, 40, 40, 40
			        4261 => x"00000000",		-- colors: 40, 40, 40, 40
			        4262 => x"00000000",		-- colors: 40, 40, 40, 40
			        4263 => x"00000000",		-- colors: 40, 40, 40, 40
			        4264 => x"00000000",		-- colors: 40, 40, 40, 40
			        4265 => x"00000000",		-- colors: 40, 40, 40, 40
			        4266 => x"00000000",		-- colors: 40, 40, 40, 40
			        4267 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4268 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4269 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4270 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4271 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4272 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4273 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4274 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4275 => x"00000000",		-- colors: 40, 40, 40, 40
			        4276 => x"00000000",		-- colors: 40, 40, 40, 40
			        4277 => x"00000000",		-- colors: 40, 40, 40, 40
			        4278 => x"00000000",		-- colors: 40, 40, 40, 40
			        4279 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4280 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4281 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4282 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4283 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4284 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4285 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4286 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60

			                --  sprite 63
			        4287 => x"00000000",		-- colors: 40, 40, 40, 40
			        4288 => x"00000000",		-- colors: 40, 40, 40, 40
			        4289 => x"00000000",		-- colors: 40, 40, 40, 40
			        4290 => x"00000000",		-- colors: 40, 40, 40, 40
			        4291 => x"00000000",		-- colors: 40, 40, 40, 40
			        4292 => x"00000000",		-- colors: 40, 40, 40, 40
			        4293 => x"00000000",		-- colors: 40, 40, 40, 40
			        4294 => x"00000000",		-- colors: 40, 40, 40, 40
			        4295 => x"00000000",		-- colors: 40, 40, 40, 40
			        4296 => x"00000000",		-- colors: 40, 40, 40, 40
			        4297 => x"00000000",		-- colors: 40, 40, 40, 40
			        4298 => x"00000000",		-- colors: 40, 40, 40, 40
			        4299 => x"00000000",		-- colors: 40, 40, 40, 40
			        4300 => x"00000000",		-- colors: 40, 40, 40, 40
			        4301 => x"00000000",		-- colors: 40, 40, 40, 40
			        4302 => x"00000000",		-- colors: 40, 40, 40, 40
			        4303 => x"00000000",		-- colors: 40, 40, 40, 40
			        4304 => x"00000000",		-- colors: 40, 40, 40, 40
			        4305 => x"00000000",		-- colors: 40, 40, 40, 40
			        4306 => x"00000000",		-- colors: 40, 40, 40, 40
			        4307 => x"00000000",		-- colors: 40, 40, 40, 40
			        4308 => x"00000000",		-- colors: 40, 40, 40, 40
			        4309 => x"00000000",		-- colors: 40, 40, 40, 40
			        4310 => x"00000000",		-- colors: 40, 40, 40, 40
			        4311 => x"00000000",		-- colors: 40, 40, 40, 40
			        4312 => x"00000000",		-- colors: 40, 40, 40, 40
			        4313 => x"00000000",		-- colors: 40, 40, 40, 40
			        4314 => x"00000000",		-- colors: 40, 40, 40, 40
			        4315 => x"00000000",		-- colors: 40, 40, 40, 40
			        4316 => x"00000000",		-- colors: 40, 40, 40, 40
			        4317 => x"00000000",		-- colors: 40, 40, 40, 40
			        4318 => x"00000000",		-- colors: 40, 40, 40, 40
			        4319 => x"00000000",		-- colors: 40, 40, 40, 40
			        4320 => x"00000000",		-- colors: 40, 40, 40, 40
			        4321 => x"00000000",		-- colors: 40, 40, 40, 40
			        4322 => x"00000000",		-- colors: 40, 40, 40, 40
			        4323 => x"00000000",		-- colors: 40, 40, 40, 40
			        4324 => x"00000000",		-- colors: 40, 40, 40, 40
			        4325 => x"00000000",		-- colors: 40, 40, 40, 40
			        4326 => x"00000000",		-- colors: 40, 40, 40, 40
			        4327 => x"00000000",		-- colors: 40, 40, 40, 40
			        4328 => x"00000000",		-- colors: 40, 40, 40, 40
			        4329 => x"00000000",		-- colors: 40, 40, 40, 40
			        4330 => x"00000000",		-- colors: 40, 40, 40, 40
			        4331 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4332 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4333 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4334 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4335 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4336 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4337 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4338 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4339 => x"00000000",		-- colors: 40, 40, 40, 40
			        4340 => x"00000000",		-- colors: 40, 40, 40, 40
			        4341 => x"00000000",		-- colors: 40, 40, 40, 40
			        4342 => x"00000000",		-- colors: 40, 40, 40, 40
			        4343 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4344 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4345 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4346 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4347 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4348 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4349 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4350 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60

			                --  sprite 64
			        4351 => x"00000000",		-- colors: 40, 40, 40, 40
			        4352 => x"00000000",		-- colors: 40, 40, 40, 40
			        4353 => x"00000000",		-- colors: 40, 40, 40, 40
			        4354 => x"00000000",		-- colors: 40, 40, 40, 40
			        4355 => x"00000000",		-- colors: 40, 40, 40, 40
			        4356 => x"00000000",		-- colors: 40, 40, 40, 40
			        4357 => x"00000000",		-- colors: 40, 40, 40, 40
			        4358 => x"00000000",		-- colors: 40, 40, 40, 40
			        4359 => x"32323232",		-- colors: 50, 50, 50, 50
			        4360 => x"32323232",		-- colors: 50, 50, 50, 50
			        4361 => x"32323232",		-- colors: 50, 50, 50, 50
			        4362 => x"32323232",		-- colors: 50, 50, 50, 50
			        4363 => x"00000000",		-- colors: 40, 40, 40, 40
			        4364 => x"00000000",		-- colors: 40, 40, 40, 40
			        4365 => x"00000000",		-- colors: 40, 40, 40, 40
			        4366 => x"00000000",		-- colors: 40, 40, 40, 40
			        4367 => x"00000000",		-- colors: 40, 40, 40, 40
			        4368 => x"00000000",		-- colors: 40, 40, 40, 40
			        4369 => x"00000000",		-- colors: 40, 40, 40, 40
			        4370 => x"00000000",		-- colors: 40, 40, 40, 40
			        4371 => x"00000000",		-- colors: 40, 40, 40, 40
			        4372 => x"00000000",		-- colors: 40, 40, 40, 40
			        4373 => x"00000000",		-- colors: 40, 40, 40, 40
			        4374 => x"00000000",		-- colors: 40, 40, 40, 40
			        4375 => x"32323232",		-- colors: 50, 50, 50, 50
			        4376 => x"32323232",		-- colors: 50, 50, 50, 50
			        4377 => x"32323232",		-- colors: 50, 50, 50, 50
			        4378 => x"32323232",		-- colors: 50, 50, 50, 50
			        4379 => x"00000000",		-- colors: 40, 40, 40, 40
			        4380 => x"00000000",		-- colors: 40, 40, 40, 40
			        4381 => x"00000000",		-- colors: 40, 40, 40, 40
			        4382 => x"00000000",		-- colors: 40, 40, 40, 40
			        4383 => x"00000000",		-- colors: 40, 40, 40, 40
			        4384 => x"00000000",		-- colors: 40, 40, 40, 40
			        4385 => x"00000000",		-- colors: 40, 40, 40, 40
			        4386 => x"00000000",		-- colors: 40, 40, 40, 40
			        4387 => x"00000000",		-- colors: 40, 40, 40, 40
			        4388 => x"00000000",		-- colors: 40, 40, 40, 40
			        4389 => x"00000000",		-- colors: 40, 40, 40, 40
			        4390 => x"00000000",		-- colors: 40, 40, 40, 40
			        4391 => x"32323232",		-- colors: 50, 50, 50, 50
			        4392 => x"32323232",		-- colors: 50, 50, 50, 50
			        4393 => x"32323232",		-- colors: 50, 50, 50, 50
			        4394 => x"32323232",		-- colors: 50, 50, 50, 50
			        4395 => x"00000000",		-- colors: 40, 40, 40, 40
			        4396 => x"00000000",		-- colors: 40, 40, 40, 40
			        4397 => x"00000000",		-- colors: 40, 40, 40, 40
			        4398 => x"00000000",		-- colors: 40, 40, 40, 40
			        4399 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4400 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4401 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4402 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4403 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4404 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4405 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4406 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4407 => x"00000000",		-- colors: 40, 40, 40, 40
			        4408 => x"00000000",		-- colors: 40, 40, 40, 40
			        4409 => x"00000000",		-- colors: 40, 40, 40, 40
			        4410 => x"00000000",		-- colors: 40, 40, 40, 40
			        4411 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4412 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4413 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4414 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60

			                --  sprite 65
			        4415 => x"00000000",		-- colors: 40, 40, 40, 40
			        4416 => x"00000000",		-- colors: 40, 40, 40, 40
			        4417 => x"00000000",		-- colors: 40, 40, 40, 40
			        4418 => x"00000000",		-- colors: 40, 40, 40, 40
			        4419 => x"00000000",		-- colors: 40, 40, 40, 40
			        4420 => x"00000000",		-- colors: 40, 40, 40, 40
			        4421 => x"00000000",		-- colors: 40, 40, 40, 40
			        4422 => x"00000000",		-- colors: 40, 40, 40, 40
			        4423 => x"00000000",		-- colors: 40, 40, 40, 40
			        4424 => x"00000000",		-- colors: 40, 40, 40, 40
			        4425 => x"00000000",		-- colors: 40, 40, 40, 40
			        4426 => x"00000000",		-- colors: 40, 40, 40, 40
			        4427 => x"00000000",		-- colors: 40, 40, 40, 40
			        4428 => x"00000000",		-- colors: 40, 40, 40, 40
			        4429 => x"00000000",		-- colors: 40, 40, 40, 40
			        4430 => x"00000000",		-- colors: 40, 40, 40, 40
			        4431 => x"00000000",		-- colors: 40, 40, 40, 40
			        4432 => x"00000000",		-- colors: 40, 40, 40, 40
			        4433 => x"00000000",		-- colors: 40, 40, 40, 40
			        4434 => x"00000000",		-- colors: 40, 40, 40, 40
			        4435 => x"00000000",		-- colors: 40, 40, 40, 40
			        4436 => x"00000000",		-- colors: 40, 40, 40, 40
			        4437 => x"00000000",		-- colors: 40, 40, 40, 40
			        4438 => x"00000000",		-- colors: 40, 40, 40, 40
			        4439 => x"00000000",		-- colors: 40, 40, 40, 40
			        4440 => x"00000000",		-- colors: 40, 40, 40, 40
			        4441 => x"00000000",		-- colors: 40, 40, 40, 40
			        4442 => x"00000000",		-- colors: 40, 40, 40, 40
			        4443 => x"00000000",		-- colors: 40, 40, 40, 40
			        4444 => x"00000000",		-- colors: 40, 40, 40, 40
			        4445 => x"00000000",		-- colors: 40, 40, 40, 40
			        4446 => x"00000000",		-- colors: 40, 40, 40, 40
			        4447 => x"00000000",		-- colors: 40, 40, 40, 40
			        4448 => x"00000000",		-- colors: 40, 40, 40, 40
			        4449 => x"00000000",		-- colors: 40, 40, 40, 40
			        4450 => x"00000000",		-- colors: 40, 40, 40, 40
			        4451 => x"00000000",		-- colors: 40, 40, 40, 40
			        4452 => x"00000000",		-- colors: 40, 40, 40, 40
			        4453 => x"00000000",		-- colors: 40, 40, 40, 40
			        4454 => x"00000000",		-- colors: 40, 40, 40, 40
			        4455 => x"00000000",		-- colors: 40, 40, 40, 40
			        4456 => x"00000000",		-- colors: 40, 40, 40, 40
			        4457 => x"00000000",		-- colors: 40, 40, 40, 40
			        4458 => x"00000000",		-- colors: 40, 40, 40, 40
			        4459 => x"00000000",		-- colors: 40, 40, 40, 40
			        4460 => x"00000000",		-- colors: 40, 40, 40, 40
			        4461 => x"00000000",		-- colors: 40, 40, 40, 40
			        4462 => x"00000000",		-- colors: 40, 40, 40, 40
			        4463 => x"00000000",		-- colors: 40, 40, 40, 40
			        4464 => x"00000000",		-- colors: 40, 40, 40, 40
			        4465 => x"00000000",		-- colors: 40, 40, 40, 40
			        4466 => x"00000000",		-- colors: 40, 40, 40, 40
			        4467 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4468 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4469 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4470 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4471 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4472 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4473 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4474 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4475 => x"00000000",		-- colors: 40, 40, 40, 40
			        4476 => x"00000000",		-- colors: 40, 40, 40, 40
			        4477 => x"00000000",		-- colors: 40, 40, 40, 40
			        4478 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 66
			        4479 => x"00000000",		-- colors: 40, 40, 40, 40
			        4480 => x"00000000",		-- colors: 40, 40, 40, 40
			        4481 => x"00000000",		-- colors: 40, 40, 40, 40
			        4482 => x"00000000",		-- colors: 40, 40, 40, 40
			        4483 => x"00000000",		-- colors: 40, 40, 40, 40
			        4484 => x"00000000",		-- colors: 40, 40, 40, 40
			        4485 => x"00000000",		-- colors: 40, 40, 40, 40
			        4486 => x"00000000",		-- colors: 40, 40, 40, 40
			        4487 => x"00000000",		-- colors: 40, 40, 40, 40
			        4488 => x"00000000",		-- colors: 40, 40, 40, 40
			        4489 => x"00000000",		-- colors: 40, 40, 40, 40
			        4490 => x"00000000",		-- colors: 40, 40, 40, 40
			        4491 => x"00000000",		-- colors: 40, 40, 40, 40
			        4492 => x"00000000",		-- colors: 40, 40, 40, 40
			        4493 => x"00000000",		-- colors: 40, 40, 40, 40
			        4494 => x"00000000",		-- colors: 40, 40, 40, 40
			        4495 => x"00000000",		-- colors: 40, 40, 40, 40
			        4496 => x"00000000",		-- colors: 40, 40, 40, 40
			        4497 => x"00000000",		-- colors: 40, 40, 40, 40
			        4498 => x"00000000",		-- colors: 40, 40, 40, 40
			        4499 => x"00000000",		-- colors: 40, 40, 40, 40
			        4500 => x"00000000",		-- colors: 40, 40, 40, 40
			        4501 => x"00000000",		-- colors: 40, 40, 40, 40
			        4502 => x"00000000",		-- colors: 40, 40, 40, 40
			        4503 => x"00000000",		-- colors: 40, 40, 40, 40
			        4504 => x"00000000",		-- colors: 40, 40, 40, 40
			        4505 => x"00000000",		-- colors: 40, 40, 40, 40
			        4506 => x"00000000",		-- colors: 40, 40, 40, 40
			        4507 => x"00000000",		-- colors: 40, 40, 40, 40
			        4508 => x"00000000",		-- colors: 40, 40, 40, 40
			        4509 => x"00000000",		-- colors: 40, 40, 40, 40
			        4510 => x"00000000",		-- colors: 40, 40, 40, 40
			        4511 => x"00000000",		-- colors: 40, 40, 40, 40
			        4512 => x"00000000",		-- colors: 40, 40, 40, 40
			        4513 => x"00000000",		-- colors: 40, 40, 40, 40
			        4514 => x"00000000",		-- colors: 40, 40, 40, 40
			        4515 => x"00000000",		-- colors: 40, 40, 40, 40
			        4516 => x"00000000",		-- colors: 40, 40, 40, 40
			        4517 => x"00000000",		-- colors: 40, 40, 40, 40
			        4518 => x"00000000",		-- colors: 40, 40, 40, 40
			        4519 => x"00000000",		-- colors: 40, 40, 40, 40
			        4520 => x"00000000",		-- colors: 40, 40, 40, 40
			        4521 => x"00000000",		-- colors: 40, 40, 40, 40
			        4522 => x"00000000",		-- colors: 40, 40, 40, 40
			        4523 => x"00000000",		-- colors: 40, 40, 40, 40
			        4524 => x"00000000",		-- colors: 40, 40, 40, 40
			        4525 => x"00000000",		-- colors: 40, 40, 40, 40
			        4526 => x"00000000",		-- colors: 40, 40, 40, 40
			        4527 => x"00000000",		-- colors: 40, 40, 40, 40
			        4528 => x"00000000",		-- colors: 40, 40, 40, 40
			        4529 => x"00000000",		-- colors: 40, 40, 40, 40
			        4530 => x"00000000",		-- colors: 40, 40, 40, 40
			        4531 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4532 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4533 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4534 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4535 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4536 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4537 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4538 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4539 => x"00000000",		-- colors: 40, 40, 40, 40
			        4540 => x"00000000",		-- colors: 40, 40, 40, 40
			        4541 => x"00000000",		-- colors: 40, 40, 40, 40
			        4542 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 67
			        4543 => x"00000000",		-- colors: 40, 40, 40, 40
			        4544 => x"00000000",		-- colors: 40, 40, 40, 40
			        4545 => x"00000000",		-- colors: 40, 40, 40, 40
			        4546 => x"00000000",		-- colors: 40, 40, 40, 40
			        4547 => x"00000000",		-- colors: 40, 40, 40, 40
			        4548 => x"00000000",		-- colors: 40, 40, 40, 40
			        4549 => x"00000000",		-- colors: 40, 40, 40, 40
			        4550 => x"00000000",		-- colors: 40, 40, 40, 40
			        4551 => x"00000000",		-- colors: 40, 40, 40, 40
			        4552 => x"00000000",		-- colors: 40, 40, 40, 40
			        4553 => x"00000000",		-- colors: 40, 40, 40, 40
			        4554 => x"00000000",		-- colors: 40, 40, 40, 40
			        4555 => x"00000000",		-- colors: 40, 40, 40, 40
			        4556 => x"00000000",		-- colors: 40, 40, 40, 40
			        4557 => x"00000000",		-- colors: 40, 40, 40, 40
			        4558 => x"00000000",		-- colors: 40, 40, 40, 40
			        4559 => x"00000000",		-- colors: 40, 40, 40, 40
			        4560 => x"00000000",		-- colors: 40, 40, 40, 40
			        4561 => x"00000000",		-- colors: 40, 40, 40, 40
			        4562 => x"00000000",		-- colors: 40, 40, 40, 40
			        4563 => x"00000000",		-- colors: 40, 40, 40, 40
			        4564 => x"00000000",		-- colors: 40, 40, 40, 40
			        4565 => x"00000000",		-- colors: 40, 40, 40, 40
			        4566 => x"00000000",		-- colors: 40, 40, 40, 40
			        4567 => x"00000000",		-- colors: 40, 40, 40, 40
			        4568 => x"00000000",		-- colors: 40, 40, 40, 40
			        4569 => x"00000000",		-- colors: 40, 40, 40, 40
			        4570 => x"00000000",		-- colors: 40, 40, 40, 40
			        4571 => x"00000000",		-- colors: 40, 40, 40, 40
			        4572 => x"00000000",		-- colors: 40, 40, 40, 40
			        4573 => x"00000000",		-- colors: 40, 40, 40, 40
			        4574 => x"00000000",		-- colors: 40, 40, 40, 40
			        4575 => x"00000000",		-- colors: 40, 40, 40, 40
			        4576 => x"00000000",		-- colors: 40, 40, 40, 40
			        4577 => x"00000000",		-- colors: 40, 40, 40, 40
			        4578 => x"00000000",		-- colors: 40, 40, 40, 40
			        4579 => x"00000000",		-- colors: 40, 40, 40, 40
			        4580 => x"00000000",		-- colors: 40, 40, 40, 40
			        4581 => x"00000000",		-- colors: 40, 40, 40, 40
			        4582 => x"00000000",		-- colors: 40, 40, 40, 40
			        4583 => x"00000000",		-- colors: 40, 40, 40, 40
			        4584 => x"00000000",		-- colors: 40, 40, 40, 40
			        4585 => x"00000000",		-- colors: 40, 40, 40, 40
			        4586 => x"00000000",		-- colors: 40, 40, 40, 40
			        4587 => x"00000000",		-- colors: 40, 40, 40, 40
			        4588 => x"00000000",		-- colors: 40, 40, 40, 40
			        4589 => x"00000000",		-- colors: 40, 40, 40, 40
			        4590 => x"00000000",		-- colors: 40, 40, 40, 40
			        4591 => x"00000000",		-- colors: 40, 40, 40, 40
			        4592 => x"00000000",		-- colors: 40, 40, 40, 40
			        4593 => x"00000000",		-- colors: 40, 40, 40, 40
			        4594 => x"00000000",		-- colors: 40, 40, 40, 40
			        4595 => x"00000000",		-- colors: 40, 40, 40, 40
			        4596 => x"00000000",		-- colors: 40, 40, 40, 40
			        4597 => x"00000000",		-- colors: 40, 40, 40, 40
			        4598 => x"00000000",		-- colors: 40, 40, 40, 40
			        4599 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4600 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4601 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4602 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4603 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4604 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4605 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4606 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60

			                --  sprite 68
			        4607 => x"00000000",		-- colors: 40, 40, 40, 40
			        4608 => x"00000000",		-- colors: 40, 40, 40, 40
			        4609 => x"00000000",		-- colors: 40, 40, 40, 40
			        4610 => x"00000000",		-- colors: 40, 40, 40, 40
			        4611 => x"00000000",		-- colors: 40, 40, 40, 40
			        4612 => x"00000000",		-- colors: 40, 40, 40, 40
			        4613 => x"00000000",		-- colors: 40, 40, 40, 40
			        4614 => x"00000000",		-- colors: 40, 40, 40, 40
			        4615 => x"00000000",		-- colors: 40, 40, 40, 40
			        4616 => x"00000000",		-- colors: 40, 40, 40, 40
			        4617 => x"00000000",		-- colors: 40, 40, 40, 40
			        4618 => x"00000000",		-- colors: 40, 40, 40, 40
			        4619 => x"00000000",		-- colors: 40, 40, 40, 40
			        4620 => x"00000000",		-- colors: 40, 40, 40, 40
			        4621 => x"00000000",		-- colors: 40, 40, 40, 40
			        4622 => x"00000000",		-- colors: 40, 40, 40, 40
			        4623 => x"00000000",		-- colors: 40, 40, 40, 40
			        4624 => x"00000000",		-- colors: 40, 40, 40, 40
			        4625 => x"00000000",		-- colors: 40, 40, 40, 40
			        4626 => x"00000000",		-- colors: 40, 40, 40, 40
			        4627 => x"00000000",		-- colors: 40, 40, 40, 40
			        4628 => x"00000000",		-- colors: 40, 40, 40, 40
			        4629 => x"00000000",		-- colors: 40, 40, 40, 40
			        4630 => x"00000000",		-- colors: 40, 40, 40, 40
			        4631 => x"00000000",		-- colors: 40, 40, 40, 40
			        4632 => x"00000000",		-- colors: 40, 40, 40, 40
			        4633 => x"00000000",		-- colors: 40, 40, 40, 40
			        4634 => x"00000000",		-- colors: 40, 40, 40, 40
			        4635 => x"00000000",		-- colors: 40, 40, 40, 40
			        4636 => x"00000000",		-- colors: 40, 40, 40, 40
			        4637 => x"00000000",		-- colors: 40, 40, 40, 40
			        4638 => x"00000000",		-- colors: 40, 40, 40, 40
			        4639 => x"00000000",		-- colors: 40, 40, 40, 40
			        4640 => x"00000000",		-- colors: 40, 40, 40, 40
			        4641 => x"00000000",		-- colors: 40, 40, 40, 40
			        4642 => x"00000000",		-- colors: 40, 40, 40, 40
			        4643 => x"00000000",		-- colors: 40, 40, 40, 40
			        4644 => x"00000000",		-- colors: 40, 40, 40, 40
			        4645 => x"00000000",		-- colors: 40, 40, 40, 40
			        4646 => x"00000000",		-- colors: 40, 40, 40, 40
			        4647 => x"00000000",		-- colors: 40, 40, 40, 40
			        4648 => x"00000000",		-- colors: 40, 40, 40, 40
			        4649 => x"00000000",		-- colors: 40, 40, 40, 40
			        4650 => x"00000000",		-- colors: 40, 40, 40, 40
			        4651 => x"00000000",		-- colors: 40, 40, 40, 40
			        4652 => x"00000000",		-- colors: 40, 40, 40, 40
			        4653 => x"00000000",		-- colors: 40, 40, 40, 40
			        4654 => x"00000000",		-- colors: 40, 40, 40, 40
			        4655 => x"00000000",		-- colors: 40, 40, 40, 40
			        4656 => x"00000000",		-- colors: 40, 40, 40, 40
			        4657 => x"00000000",		-- colors: 40, 40, 40, 40
			        4658 => x"00000000",		-- colors: 40, 40, 40, 40
			        4659 => x"00000000",		-- colors: 40, 40, 40, 40
			        4660 => x"00000000",		-- colors: 40, 40, 40, 40
			        4661 => x"00000000",		-- colors: 40, 40, 40, 40
			        4662 => x"00000000",		-- colors: 40, 40, 40, 40
			        4663 => x"00000000",		-- colors: 40, 40, 40, 40
			        4664 => x"00000000",		-- colors: 40, 40, 40, 40
			        4665 => x"00000000",		-- colors: 40, 40, 40, 40
			        4666 => x"00000000",		-- colors: 40, 40, 40, 40
			        4667 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4668 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4669 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4670 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60

			                --  sprite 69
			        4671 => x"00000000",		-- colors: 40, 40, 40, 40
			        4672 => x"00000000",		-- colors: 40, 40, 40, 40
			        4673 => x"00000000",		-- colors: 40, 40, 40, 40
			        4674 => x"00000000",		-- colors: 40, 40, 40, 40
			        4675 => x"00000000",		-- colors: 40, 40, 40, 40
			        4676 => x"00000000",		-- colors: 40, 40, 40, 40
			        4677 => x"00000000",		-- colors: 40, 40, 40, 40
			        4678 => x"00000000",		-- colors: 40, 40, 40, 40
			        4679 => x"00000000",		-- colors: 40, 40, 40, 40
			        4680 => x"00000000",		-- colors: 40, 40, 40, 40
			        4681 => x"00000000",		-- colors: 40, 40, 40, 40
			        4682 => x"00000000",		-- colors: 40, 40, 40, 40
			        4683 => x"00000000",		-- colors: 40, 40, 40, 40
			        4684 => x"00000000",		-- colors: 40, 40, 40, 40
			        4685 => x"00000000",		-- colors: 40, 40, 40, 40
			        4686 => x"00000000",		-- colors: 40, 40, 40, 40
			        4687 => x"00000000",		-- colors: 40, 40, 40, 40
			        4688 => x"00000000",		-- colors: 40, 40, 40, 40
			        4689 => x"00000000",		-- colors: 40, 40, 40, 40
			        4690 => x"00000000",		-- colors: 40, 40, 40, 40
			        4691 => x"00000000",		-- colors: 40, 40, 40, 40
			        4692 => x"00000000",		-- colors: 40, 40, 40, 40
			        4693 => x"00000000",		-- colors: 40, 40, 40, 40
			        4694 => x"00000000",		-- colors: 40, 40, 40, 40
			        4695 => x"00000000",		-- colors: 40, 40, 40, 40
			        4696 => x"00000000",		-- colors: 40, 40, 40, 40
			        4697 => x"00000000",		-- colors: 40, 40, 40, 40
			        4698 => x"00000000",		-- colors: 40, 40, 40, 40
			        4699 => x"00000000",		-- colors: 40, 40, 40, 40
			        4700 => x"00000000",		-- colors: 40, 40, 40, 40
			        4701 => x"00000000",		-- colors: 40, 40, 40, 40
			        4702 => x"00000000",		-- colors: 40, 40, 40, 40
			        4703 => x"00000000",		-- colors: 40, 40, 40, 40
			        4704 => x"00000000",		-- colors: 40, 40, 40, 40
			        4705 => x"00000000",		-- colors: 40, 40, 40, 40
			        4706 => x"00000000",		-- colors: 40, 40, 40, 40
			        4707 => x"00000000",		-- colors: 40, 40, 40, 40
			        4708 => x"00000000",		-- colors: 40, 40, 40, 40
			        4709 => x"00000000",		-- colors: 40, 40, 40, 40
			        4710 => x"00000000",		-- colors: 40, 40, 40, 40
			        4711 => x"00000000",		-- colors: 40, 40, 40, 40
			        4712 => x"00000000",		-- colors: 40, 40, 40, 40
			        4713 => x"00000000",		-- colors: 40, 40, 40, 40
			        4714 => x"00000000",		-- colors: 40, 40, 40, 40
			        4715 => x"00000000",		-- colors: 40, 40, 40, 40
			        4716 => x"00000000",		-- colors: 40, 40, 40, 40
			        4717 => x"00000000",		-- colors: 40, 40, 40, 40
			        4718 => x"00000000",		-- colors: 40, 40, 40, 40
			        4719 => x"00000000",		-- colors: 40, 40, 40, 40
			        4720 => x"00000000",		-- colors: 40, 40, 40, 40
			        4721 => x"00000000",		-- colors: 40, 40, 40, 40
			        4722 => x"00000000",		-- colors: 40, 40, 40, 40
			        4723 => x"00000000",		-- colors: 40, 40, 40, 40
			        4724 => x"00000000",		-- colors: 40, 40, 40, 40
			        4725 => x"00000000",		-- colors: 40, 40, 40, 40
			        4726 => x"00000000",		-- colors: 40, 40, 40, 40
			        4727 => x"00000000",		-- colors: 40, 40, 40, 40
			        4728 => x"00000000",		-- colors: 40, 40, 40, 40
			        4729 => x"00000000",		-- colors: 40, 40, 40, 40
			        4730 => x"00000000",		-- colors: 40, 40, 40, 40
			        4731 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4732 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4733 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4734 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60

			                --  sprite 70
			        4735 => x"00000000",		-- colors: 40, 40, 40, 40
			        4736 => x"00000000",		-- colors: 40, 40, 40, 40
			        4737 => x"00000000",		-- colors: 40, 40, 40, 40
			        4738 => x"00000000",		-- colors: 40, 40, 40, 40
			        4739 => x"00000000",		-- colors: 40, 40, 40, 40
			        4740 => x"00000000",		-- colors: 40, 40, 40, 40
			        4741 => x"00000000",		-- colors: 40, 40, 40, 40
			        4742 => x"00000000",		-- colors: 40, 40, 40, 40
			        4743 => x"00000000",		-- colors: 40, 40, 40, 40
			        4744 => x"00000000",		-- colors: 40, 40, 40, 40
			        4745 => x"00000000",		-- colors: 40, 40, 40, 40
			        4746 => x"00000000",		-- colors: 40, 40, 40, 40
			        4747 => x"00000000",		-- colors: 40, 40, 40, 40
			        4748 => x"00000000",		-- colors: 40, 40, 40, 40
			        4749 => x"00000000",		-- colors: 40, 40, 40, 40
			        4750 => x"00000000",		-- colors: 40, 40, 40, 40
			        4751 => x"00000000",		-- colors: 40, 40, 40, 40
			        4752 => x"00000000",		-- colors: 40, 40, 40, 40
			        4753 => x"00000000",		-- colors: 40, 40, 40, 40
			        4754 => x"00000000",		-- colors: 40, 40, 40, 40
			        4755 => x"00000000",		-- colors: 40, 40, 40, 40
			        4756 => x"00000000",		-- colors: 40, 40, 40, 40
			        4757 => x"00000000",		-- colors: 40, 40, 40, 40
			        4758 => x"00000000",		-- colors: 40, 40, 40, 40
			        4759 => x"00000000",		-- colors: 40, 40, 40, 40
			        4760 => x"00000000",		-- colors: 40, 40, 40, 40
			        4761 => x"00000000",		-- colors: 40, 40, 40, 40
			        4762 => x"00000000",		-- colors: 40, 40, 40, 40
			        4763 => x"00000000",		-- colors: 40, 40, 40, 40
			        4764 => x"00000000",		-- colors: 40, 40, 40, 40
			        4765 => x"00000000",		-- colors: 40, 40, 40, 40
			        4766 => x"00000000",		-- colors: 40, 40, 40, 40
			        4767 => x"00000000",		-- colors: 40, 40, 40, 40
			        4768 => x"00000000",		-- colors: 40, 40, 40, 40
			        4769 => x"00000000",		-- colors: 40, 40, 40, 40
			        4770 => x"00000000",		-- colors: 40, 40, 40, 40
			        4771 => x"00000000",		-- colors: 40, 40, 40, 40
			        4772 => x"00000000",		-- colors: 40, 40, 40, 40
			        4773 => x"00000000",		-- colors: 40, 40, 40, 40
			        4774 => x"00000000",		-- colors: 40, 40, 40, 40
			        4775 => x"32323232",		-- colors: 50, 50, 50, 50
			        4776 => x"32323232",		-- colors: 50, 50, 50, 50
			        4777 => x"32323232",		-- colors: 50, 50, 50, 50
			        4778 => x"32323232",		-- colors: 50, 50, 50, 50
			        4779 => x"00000000",		-- colors: 40, 40, 40, 40
			        4780 => x"00000000",		-- colors: 40, 40, 40, 40
			        4781 => x"00000000",		-- colors: 40, 40, 40, 40
			        4782 => x"00000000",		-- colors: 40, 40, 40, 40
			        4783 => x"00000000",		-- colors: 40, 40, 40, 40
			        4784 => x"00000000",		-- colors: 40, 40, 40, 40
			        4785 => x"00000000",		-- colors: 40, 40, 40, 40
			        4786 => x"00000000",		-- colors: 40, 40, 40, 40
			        4787 => x"00000000",		-- colors: 40, 40, 40, 40
			        4788 => x"00000000",		-- colors: 40, 40, 40, 40
			        4789 => x"00000000",		-- colors: 40, 40, 40, 40
			        4790 => x"00000000",		-- colors: 40, 40, 40, 40
			        4791 => x"32323232",		-- colors: 50, 50, 50, 50
			        4792 => x"32323232",		-- colors: 50, 50, 50, 50
			        4793 => x"32323232",		-- colors: 50, 50, 50, 50
			        4794 => x"32323232",		-- colors: 50, 50, 50, 50
			        4795 => x"00000000",		-- colors: 40, 40, 40, 40
			        4796 => x"00000000",		-- colors: 40, 40, 40, 40
			        4797 => x"00000000",		-- colors: 40, 40, 40, 40
			        4798 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 71
			        4799 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4800 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4801 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4802 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4803 => x"00000000",		-- colors: 40, 40, 40, 40
			        4804 => x"00000000",		-- colors: 40, 40, 40, 40
			        4805 => x"00000000",		-- colors: 40, 40, 40, 40
			        4806 => x"00000000",		-- colors: 40, 40, 40, 40
			        4807 => x"00000000",		-- colors: 40, 40, 40, 40
			        4808 => x"00000000",		-- colors: 40, 40, 40, 40
			        4809 => x"00000000",		-- colors: 40, 40, 40, 40
			        4810 => x"00000000",		-- colors: 40, 40, 40, 40
			        4811 => x"00000000",		-- colors: 40, 40, 40, 40
			        4812 => x"00000000",		-- colors: 40, 40, 40, 40
			        4813 => x"00000000",		-- colors: 40, 40, 40, 40
			        4814 => x"00000000",		-- colors: 40, 40, 40, 40
			        4815 => x"00000000",		-- colors: 40, 40, 40, 40
			        4816 => x"00000000",		-- colors: 40, 40, 40, 40
			        4817 => x"00000000",		-- colors: 40, 40, 40, 40
			        4818 => x"00000000",		-- colors: 40, 40, 40, 40
			        4819 => x"00000000",		-- colors: 40, 40, 40, 40
			        4820 => x"00000000",		-- colors: 40, 40, 40, 40
			        4821 => x"00000000",		-- colors: 40, 40, 40, 40
			        4822 => x"00000000",		-- colors: 40, 40, 40, 40
			        4823 => x"00000000",		-- colors: 40, 40, 40, 40
			        4824 => x"00000000",		-- colors: 40, 40, 40, 40
			        4825 => x"00000000",		-- colors: 40, 40, 40, 40
			        4826 => x"00000000",		-- colors: 40, 40, 40, 40
			        4827 => x"00000000",		-- colors: 40, 40, 40, 40
			        4828 => x"00000000",		-- colors: 40, 40, 40, 40
			        4829 => x"00000000",		-- colors: 40, 40, 40, 40
			        4830 => x"00000000",		-- colors: 40, 40, 40, 40
			        4831 => x"00000000",		-- colors: 40, 40, 40, 40
			        4832 => x"00000000",		-- colors: 40, 40, 40, 40
			        4833 => x"00000000",		-- colors: 40, 40, 40, 40
			        4834 => x"00000000",		-- colors: 40, 40, 40, 40
			        4835 => x"00000000",		-- colors: 40, 40, 40, 40
			        4836 => x"00000000",		-- colors: 40, 40, 40, 40
			        4837 => x"00000000",		-- colors: 40, 40, 40, 40
			        4838 => x"00000000",		-- colors: 40, 40, 40, 40
			        4839 => x"00000000",		-- colors: 40, 40, 40, 40
			        4840 => x"00000000",		-- colors: 40, 40, 40, 40
			        4841 => x"00000000",		-- colors: 40, 40, 40, 40
			        4842 => x"00000000",		-- colors: 40, 40, 40, 40
			        4843 => x"00000000",		-- colors: 40, 40, 40, 40
			        4844 => x"00000000",		-- colors: 40, 40, 40, 40
			        4845 => x"00000000",		-- colors: 40, 40, 40, 40
			        4846 => x"00000000",		-- colors: 40, 40, 40, 40
			        4847 => x"00000000",		-- colors: 40, 40, 40, 40
			        4848 => x"00000000",		-- colors: 40, 40, 40, 40
			        4849 => x"00000000",		-- colors: 40, 40, 40, 40
			        4850 => x"00000000",		-- colors: 40, 40, 40, 40
			        4851 => x"00000000",		-- colors: 40, 40, 40, 40
			        4852 => x"00000000",		-- colors: 40, 40, 40, 40
			        4853 => x"00000000",		-- colors: 40, 40, 40, 40
			        4854 => x"00000000",		-- colors: 40, 40, 40, 40
			        4855 => x"00000000",		-- colors: 40, 40, 40, 40
			        4856 => x"00000000",		-- colors: 40, 40, 40, 40
			        4857 => x"00000000",		-- colors: 40, 40, 40, 40
			        4858 => x"00000000",		-- colors: 40, 40, 40, 40
			        4859 => x"00000000",		-- colors: 40, 40, 40, 40
			        4860 => x"00000000",		-- colors: 40, 40, 40, 40
			        4861 => x"00000000",		-- colors: 40, 40, 40, 40
			        4862 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 72
			        4863 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4864 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4865 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4866 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4867 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4868 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4869 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4870 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4871 => x"00000000",		-- colors: 40, 40, 40, 40
			        4872 => x"00000000",		-- colors: 40, 40, 40, 40
			        4873 => x"00000000",		-- colors: 40, 40, 40, 40
			        4874 => x"00000000",		-- colors: 40, 40, 40, 40
			        4875 => x"00000000",		-- colors: 40, 40, 40, 40
			        4876 => x"00000000",		-- colors: 40, 40, 40, 40
			        4877 => x"00000000",		-- colors: 40, 40, 40, 40
			        4878 => x"00000000",		-- colors: 40, 40, 40, 40
			        4879 => x"00000000",		-- colors: 40, 40, 40, 40
			        4880 => x"00000000",		-- colors: 40, 40, 40, 40
			        4881 => x"00000000",		-- colors: 40, 40, 40, 40
			        4882 => x"00000000",		-- colors: 40, 40, 40, 40
			        4883 => x"00000000",		-- colors: 40, 40, 40, 40
			        4884 => x"00000000",		-- colors: 40, 40, 40, 40
			        4885 => x"00000000",		-- colors: 40, 40, 40, 40
			        4886 => x"00000000",		-- colors: 40, 40, 40, 40
			        4887 => x"00000000",		-- colors: 40, 40, 40, 40
			        4888 => x"00000000",		-- colors: 40, 40, 40, 40
			        4889 => x"00000000",		-- colors: 40, 40, 40, 40
			        4890 => x"00000000",		-- colors: 40, 40, 40, 40
			        4891 => x"00000000",		-- colors: 40, 40, 40, 40
			        4892 => x"00000000",		-- colors: 40, 40, 40, 40
			        4893 => x"00000000",		-- colors: 40, 40, 40, 40
			        4894 => x"00000000",		-- colors: 40, 40, 40, 40
			        4895 => x"00000000",		-- colors: 40, 40, 40, 40
			        4896 => x"00000000",		-- colors: 40, 40, 40, 40
			        4897 => x"00000000",		-- colors: 40, 40, 40, 40
			        4898 => x"00000000",		-- colors: 40, 40, 40, 40
			        4899 => x"00000000",		-- colors: 40, 40, 40, 40
			        4900 => x"00000000",		-- colors: 40, 40, 40, 40
			        4901 => x"00000000",		-- colors: 40, 40, 40, 40
			        4902 => x"00000000",		-- colors: 40, 40, 40, 40
			        4903 => x"00000000",		-- colors: 40, 40, 40, 40
			        4904 => x"00000000",		-- colors: 40, 40, 40, 40
			        4905 => x"00000000",		-- colors: 40, 40, 40, 40
			        4906 => x"00000000",		-- colors: 40, 40, 40, 40
			        4907 => x"00000000",		-- colors: 40, 40, 40, 40
			        4908 => x"00000000",		-- colors: 40, 40, 40, 40
			        4909 => x"00000000",		-- colors: 40, 40, 40, 40
			        4910 => x"00000000",		-- colors: 40, 40, 40, 40
			        4911 => x"00000000",		-- colors: 40, 40, 40, 40
			        4912 => x"00000000",		-- colors: 40, 40, 40, 40
			        4913 => x"00000000",		-- colors: 40, 40, 40, 40
			        4914 => x"00000000",		-- colors: 40, 40, 40, 40
			        4915 => x"00000000",		-- colors: 40, 40, 40, 40
			        4916 => x"00000000",		-- colors: 40, 40, 40, 40
			        4917 => x"00000000",		-- colors: 40, 40, 40, 40
			        4918 => x"00000000",		-- colors: 40, 40, 40, 40
			        4919 => x"00000000",		-- colors: 40, 40, 40, 40
			        4920 => x"00000000",		-- colors: 40, 40, 40, 40
			        4921 => x"00000000",		-- colors: 40, 40, 40, 40
			        4922 => x"00000000",		-- colors: 40, 40, 40, 40
			        4923 => x"00000000",		-- colors: 40, 40, 40, 40
			        4924 => x"00000000",		-- colors: 40, 40, 40, 40
			        4925 => x"00000000",		-- colors: 40, 40, 40, 40
			        4926 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 73
			        4927 => x"00000000",		-- colors: 40, 40, 40, 40
			        4928 => x"00000000",		-- colors: 40, 40, 40, 40
			        4929 => x"00000000",		-- colors: 40, 40, 40, 40
			        4930 => x"00000000",		-- colors: 40, 40, 40, 40
			        4931 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4932 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4933 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4934 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4935 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4936 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4937 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4938 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4939 => x"00000000",		-- colors: 40, 40, 40, 40
			        4940 => x"00000000",		-- colors: 40, 40, 40, 40
			        4941 => x"00000000",		-- colors: 40, 40, 40, 40
			        4942 => x"00000000",		-- colors: 40, 40, 40, 40
			        4943 => x"00000000",		-- colors: 40, 40, 40, 40
			        4944 => x"00000000",		-- colors: 40, 40, 40, 40
			        4945 => x"00000000",		-- colors: 40, 40, 40, 40
			        4946 => x"00000000",		-- colors: 40, 40, 40, 40
			        4947 => x"00000000",		-- colors: 40, 40, 40, 40
			        4948 => x"00000000",		-- colors: 40, 40, 40, 40
			        4949 => x"00000000",		-- colors: 40, 40, 40, 40
			        4950 => x"00000000",		-- colors: 40, 40, 40, 40
			        4951 => x"00000000",		-- colors: 40, 40, 40, 40
			        4952 => x"00000000",		-- colors: 40, 40, 40, 40
			        4953 => x"00000000",		-- colors: 40, 40, 40, 40
			        4954 => x"00000000",		-- colors: 40, 40, 40, 40
			        4955 => x"00000000",		-- colors: 40, 40, 40, 40
			        4956 => x"00000000",		-- colors: 40, 40, 40, 40
			        4957 => x"00000000",		-- colors: 40, 40, 40, 40
			        4958 => x"00000000",		-- colors: 40, 40, 40, 40
			        4959 => x"00000000",		-- colors: 40, 40, 40, 40
			        4960 => x"00000000",		-- colors: 40, 40, 40, 40
			        4961 => x"00000000",		-- colors: 40, 40, 40, 40
			        4962 => x"00000000",		-- colors: 40, 40, 40, 40
			        4963 => x"00000000",		-- colors: 40, 40, 40, 40
			        4964 => x"00000000",		-- colors: 40, 40, 40, 40
			        4965 => x"00000000",		-- colors: 40, 40, 40, 40
			        4966 => x"00000000",		-- colors: 40, 40, 40, 40
			        4967 => x"00000000",		-- colors: 40, 40, 40, 40
			        4968 => x"00000000",		-- colors: 40, 40, 40, 40
			        4969 => x"00000000",		-- colors: 40, 40, 40, 40
			        4970 => x"00000000",		-- colors: 40, 40, 40, 40
			        4971 => x"00000000",		-- colors: 40, 40, 40, 40
			        4972 => x"00000000",		-- colors: 40, 40, 40, 40
			        4973 => x"00000000",		-- colors: 40, 40, 40, 40
			        4974 => x"00000000",		-- colors: 40, 40, 40, 40
			        4975 => x"00000000",		-- colors: 40, 40, 40, 40
			        4976 => x"00000000",		-- colors: 40, 40, 40, 40
			        4977 => x"00000000",		-- colors: 40, 40, 40, 40
			        4978 => x"00000000",		-- colors: 40, 40, 40, 40
			        4979 => x"00000000",		-- colors: 40, 40, 40, 40
			        4980 => x"00000000",		-- colors: 40, 40, 40, 40
			        4981 => x"00000000",		-- colors: 40, 40, 40, 40
			        4982 => x"00000000",		-- colors: 40, 40, 40, 40
			        4983 => x"00000000",		-- colors: 40, 40, 40, 40
			        4984 => x"00000000",		-- colors: 40, 40, 40, 40
			        4985 => x"00000000",		-- colors: 40, 40, 40, 40
			        4986 => x"00000000",		-- colors: 40, 40, 40, 40
			        4987 => x"00000000",		-- colors: 40, 40, 40, 40
			        4988 => x"00000000",		-- colors: 40, 40, 40, 40
			        4989 => x"00000000",		-- colors: 40, 40, 40, 40
			        4990 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 74
			        4991 => x"00000000",		-- colors: 40, 40, 40, 40
			        4992 => x"00000000",		-- colors: 40, 40, 40, 40
			        4993 => x"00000000",		-- colors: 40, 40, 40, 40
			        4994 => x"00000000",		-- colors: 40, 40, 40, 40
			        4995 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4996 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4997 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4998 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        4999 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5000 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5001 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5002 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5003 => x"00000000",		-- colors: 40, 40, 40, 40
			        5004 => x"00000000",		-- colors: 40, 40, 40, 40
			        5005 => x"00000000",		-- colors: 40, 40, 40, 40
			        5006 => x"00000000",		-- colors: 40, 40, 40, 40
			        5007 => x"00000000",		-- colors: 40, 40, 40, 40
			        5008 => x"00000000",		-- colors: 40, 40, 40, 40
			        5009 => x"00000000",		-- colors: 40, 40, 40, 40
			        5010 => x"00000000",		-- colors: 40, 40, 40, 40
			        5011 => x"00000000",		-- colors: 40, 40, 40, 40
			        5012 => x"00000000",		-- colors: 40, 40, 40, 40
			        5013 => x"00000000",		-- colors: 40, 40, 40, 40
			        5014 => x"00000000",		-- colors: 40, 40, 40, 40
			        5015 => x"00000000",		-- colors: 40, 40, 40, 40
			        5016 => x"00000000",		-- colors: 40, 40, 40, 40
			        5017 => x"00000000",		-- colors: 40, 40, 40, 40
			        5018 => x"00000000",		-- colors: 40, 40, 40, 40
			        5019 => x"00000000",		-- colors: 40, 40, 40, 40
			        5020 => x"00000000",		-- colors: 40, 40, 40, 40
			        5021 => x"00000000",		-- colors: 40, 40, 40, 40
			        5022 => x"00000000",		-- colors: 40, 40, 40, 40
			        5023 => x"00000000",		-- colors: 40, 40, 40, 40
			        5024 => x"00000000",		-- colors: 40, 40, 40, 40
			        5025 => x"00000000",		-- colors: 40, 40, 40, 40
			        5026 => x"00000000",		-- colors: 40, 40, 40, 40
			        5027 => x"00000000",		-- colors: 40, 40, 40, 40
			        5028 => x"00000000",		-- colors: 40, 40, 40, 40
			        5029 => x"00000000",		-- colors: 40, 40, 40, 40
			        5030 => x"00000000",		-- colors: 40, 40, 40, 40
			        5031 => x"00000000",		-- colors: 40, 40, 40, 40
			        5032 => x"00000000",		-- colors: 40, 40, 40, 40
			        5033 => x"00000000",		-- colors: 40, 40, 40, 40
			        5034 => x"00000000",		-- colors: 40, 40, 40, 40
			        5035 => x"00000000",		-- colors: 40, 40, 40, 40
			        5036 => x"00000000",		-- colors: 40, 40, 40, 40
			        5037 => x"00000000",		-- colors: 40, 40, 40, 40
			        5038 => x"00000000",		-- colors: 40, 40, 40, 40
			        5039 => x"00000000",		-- colors: 40, 40, 40, 40
			        5040 => x"00000000",		-- colors: 40, 40, 40, 40
			        5041 => x"00000000",		-- colors: 40, 40, 40, 40
			        5042 => x"00000000",		-- colors: 40, 40, 40, 40
			        5043 => x"00000000",		-- colors: 40, 40, 40, 40
			        5044 => x"00000000",		-- colors: 40, 40, 40, 40
			        5045 => x"00000000",		-- colors: 40, 40, 40, 40
			        5046 => x"00000000",		-- colors: 40, 40, 40, 40
			        5047 => x"00000000",		-- colors: 40, 40, 40, 40
			        5048 => x"00000000",		-- colors: 40, 40, 40, 40
			        5049 => x"00000000",		-- colors: 40, 40, 40, 40
			        5050 => x"00000000",		-- colors: 40, 40, 40, 40
			        5051 => x"00000000",		-- colors: 40, 40, 40, 40
			        5052 => x"00000000",		-- colors: 40, 40, 40, 40
			        5053 => x"00000000",		-- colors: 40, 40, 40, 40
			        5054 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 75
			        5055 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5056 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5057 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5058 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5059 => x"00000000",		-- colors: 40, 40, 40, 40
			        5060 => x"00000000",		-- colors: 40, 40, 40, 40
			        5061 => x"00000000",		-- colors: 40, 40, 40, 40
			        5062 => x"00000000",		-- colors: 40, 40, 40, 40
			        5063 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5064 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5065 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5066 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5067 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5068 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5069 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5070 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5071 => x"00000000",		-- colors: 40, 40, 40, 40
			        5072 => x"00000000",		-- colors: 40, 40, 40, 40
			        5073 => x"00000000",		-- colors: 40, 40, 40, 40
			        5074 => x"00000000",		-- colors: 40, 40, 40, 40
			        5075 => x"00000000",		-- colors: 40, 40, 40, 40
			        5076 => x"00000000",		-- colors: 40, 40, 40, 40
			        5077 => x"00000000",		-- colors: 40, 40, 40, 40
			        5078 => x"00000000",		-- colors: 40, 40, 40, 40
			        5079 => x"00000000",		-- colors: 40, 40, 40, 40
			        5080 => x"00000000",		-- colors: 40, 40, 40, 40
			        5081 => x"00000000",		-- colors: 40, 40, 40, 40
			        5082 => x"00000000",		-- colors: 40, 40, 40, 40
			        5083 => x"00000000",		-- colors: 40, 40, 40, 40
			        5084 => x"00000000",		-- colors: 40, 40, 40, 40
			        5085 => x"00000000",		-- colors: 40, 40, 40, 40
			        5086 => x"00000000",		-- colors: 40, 40, 40, 40
			        5087 => x"00000000",		-- colors: 40, 40, 40, 40
			        5088 => x"00000000",		-- colors: 40, 40, 40, 40
			        5089 => x"00000000",		-- colors: 40, 40, 40, 40
			        5090 => x"00000000",		-- colors: 40, 40, 40, 40
			        5091 => x"00000000",		-- colors: 40, 40, 40, 40
			        5092 => x"00000000",		-- colors: 40, 40, 40, 40
			        5093 => x"00000000",		-- colors: 40, 40, 40, 40
			        5094 => x"00000000",		-- colors: 40, 40, 40, 40
			        5095 => x"00000000",		-- colors: 40, 40, 40, 40
			        5096 => x"00000000",		-- colors: 40, 40, 40, 40
			        5097 => x"00000000",		-- colors: 40, 40, 40, 40
			        5098 => x"00000000",		-- colors: 40, 40, 40, 40
			        5099 => x"00000000",		-- colors: 40, 40, 40, 40
			        5100 => x"00000000",		-- colors: 40, 40, 40, 40
			        5101 => x"00000000",		-- colors: 40, 40, 40, 40
			        5102 => x"00000000",		-- colors: 40, 40, 40, 40
			        5103 => x"00000000",		-- colors: 40, 40, 40, 40
			        5104 => x"00000000",		-- colors: 40, 40, 40, 40
			        5105 => x"00000000",		-- colors: 40, 40, 40, 40
			        5106 => x"00000000",		-- colors: 40, 40, 40, 40
			        5107 => x"00000000",		-- colors: 40, 40, 40, 40
			        5108 => x"00000000",		-- colors: 40, 40, 40, 40
			        5109 => x"00000000",		-- colors: 40, 40, 40, 40
			        5110 => x"00000000",		-- colors: 40, 40, 40, 40
			        5111 => x"00000000",		-- colors: 40, 40, 40, 40
			        5112 => x"00000000",		-- colors: 40, 40, 40, 40
			        5113 => x"00000000",		-- colors: 40, 40, 40, 40
			        5114 => x"00000000",		-- colors: 40, 40, 40, 40
			        5115 => x"00000000",		-- colors: 40, 40, 40, 40
			        5116 => x"00000000",		-- colors: 40, 40, 40, 40
			        5117 => x"00000000",		-- colors: 40, 40, 40, 40
			        5118 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 76
			        5119 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5120 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5121 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5122 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5123 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5124 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5125 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5126 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5127 => x"00000000",		-- colors: 40, 40, 40, 40
			        5128 => x"00000000",		-- colors: 40, 40, 40, 40
			        5129 => x"00000000",		-- colors: 40, 40, 40, 40
			        5130 => x"00000000",		-- colors: 40, 40, 40, 40
			        5131 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5132 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5133 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5134 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5135 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5136 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5137 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5138 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5139 => x"00000000",		-- colors: 40, 40, 40, 40
			        5140 => x"00000000",		-- colors: 40, 40, 40, 40
			        5141 => x"00000000",		-- colors: 40, 40, 40, 40
			        5142 => x"00000000",		-- colors: 40, 40, 40, 40
			        5143 => x"00000000",		-- colors: 40, 40, 40, 40
			        5144 => x"00000000",		-- colors: 40, 40, 40, 40
			        5145 => x"00000000",		-- colors: 40, 40, 40, 40
			        5146 => x"00000000",		-- colors: 40, 40, 40, 40
			        5147 => x"00000000",		-- colors: 40, 40, 40, 40
			        5148 => x"00000000",		-- colors: 40, 40, 40, 40
			        5149 => x"00000000",		-- colors: 40, 40, 40, 40
			        5150 => x"00000000",		-- colors: 40, 40, 40, 40
			        5151 => x"00000000",		-- colors: 40, 40, 40, 40
			        5152 => x"00000000",		-- colors: 40, 40, 40, 40
			        5153 => x"00000000",		-- colors: 40, 40, 40, 40
			        5154 => x"00000000",		-- colors: 40, 40, 40, 40
			        5155 => x"00000000",		-- colors: 40, 40, 40, 40
			        5156 => x"00000000",		-- colors: 40, 40, 40, 40
			        5157 => x"00000000",		-- colors: 40, 40, 40, 40
			        5158 => x"00000000",		-- colors: 40, 40, 40, 40
			        5159 => x"00000000",		-- colors: 40, 40, 40, 40
			        5160 => x"00000000",		-- colors: 40, 40, 40, 40
			        5161 => x"00000000",		-- colors: 40, 40, 40, 40
			        5162 => x"00000000",		-- colors: 40, 40, 40, 40
			        5163 => x"00000000",		-- colors: 40, 40, 40, 40
			        5164 => x"00000000",		-- colors: 40, 40, 40, 40
			        5165 => x"00000000",		-- colors: 40, 40, 40, 40
			        5166 => x"00000000",		-- colors: 40, 40, 40, 40
			        5167 => x"00000000",		-- colors: 40, 40, 40, 40
			        5168 => x"00000000",		-- colors: 40, 40, 40, 40
			        5169 => x"00000000",		-- colors: 40, 40, 40, 40
			        5170 => x"00000000",		-- colors: 40, 40, 40, 40
			        5171 => x"00000000",		-- colors: 40, 40, 40, 40
			        5172 => x"00000000",		-- colors: 40, 40, 40, 40
			        5173 => x"00000000",		-- colors: 40, 40, 40, 40
			        5174 => x"00000000",		-- colors: 40, 40, 40, 40
			        5175 => x"00000000",		-- colors: 40, 40, 40, 40
			        5176 => x"00000000",		-- colors: 40, 40, 40, 40
			        5177 => x"00000000",		-- colors: 40, 40, 40, 40
			        5178 => x"00000000",		-- colors: 40, 40, 40, 40
			        5179 => x"00000000",		-- colors: 40, 40, 40, 40
			        5180 => x"00000000",		-- colors: 40, 40, 40, 40
			        5181 => x"00000000",		-- colors: 40, 40, 40, 40
			        5182 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 77
			        5183 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5184 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5185 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5186 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5187 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5188 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5189 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5190 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5191 => x"00000000",		-- colors: 40, 40, 40, 40
			        5192 => x"00000000",		-- colors: 40, 40, 40, 40
			        5193 => x"00000000",		-- colors: 40, 40, 40, 40
			        5194 => x"00000000",		-- colors: 40, 40, 40, 40
			        5195 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5196 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5197 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5198 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5199 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5200 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5201 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5202 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5203 => x"00000000",		-- colors: 40, 40, 40, 40
			        5204 => x"00000000",		-- colors: 40, 40, 40, 40
			        5205 => x"00000000",		-- colors: 40, 40, 40, 40
			        5206 => x"00000000",		-- colors: 40, 40, 40, 40
			        5207 => x"00000000",		-- colors: 40, 40, 40, 40
			        5208 => x"00000000",		-- colors: 40, 40, 40, 40
			        5209 => x"00000000",		-- colors: 40, 40, 40, 40
			        5210 => x"00000000",		-- colors: 40, 40, 40, 40
			        5211 => x"00000000",		-- colors: 40, 40, 40, 40
			        5212 => x"00000000",		-- colors: 40, 40, 40, 40
			        5213 => x"00000000",		-- colors: 40, 40, 40, 40
			        5214 => x"00000000",		-- colors: 40, 40, 40, 40
			        5215 => x"00000000",		-- colors: 40, 40, 40, 40
			        5216 => x"00000000",		-- colors: 40, 40, 40, 40
			        5217 => x"00000000",		-- colors: 40, 40, 40, 40
			        5218 => x"00000000",		-- colors: 40, 40, 40, 40
			        5219 => x"00000000",		-- colors: 40, 40, 40, 40
			        5220 => x"00000000",		-- colors: 40, 40, 40, 40
			        5221 => x"00000000",		-- colors: 40, 40, 40, 40
			        5222 => x"00000000",		-- colors: 40, 40, 40, 40
			        5223 => x"00000000",		-- colors: 40, 40, 40, 40
			        5224 => x"00000000",		-- colors: 40, 40, 40, 40
			        5225 => x"00000000",		-- colors: 40, 40, 40, 40
			        5226 => x"00000000",		-- colors: 40, 40, 40, 40
			        5227 => x"00000000",		-- colors: 40, 40, 40, 40
			        5228 => x"00000000",		-- colors: 40, 40, 40, 40
			        5229 => x"00000000",		-- colors: 40, 40, 40, 40
			        5230 => x"00000000",		-- colors: 40, 40, 40, 40
			        5231 => x"00000000",		-- colors: 40, 40, 40, 40
			        5232 => x"00000000",		-- colors: 40, 40, 40, 40
			        5233 => x"00000000",		-- colors: 40, 40, 40, 40
			        5234 => x"00000000",		-- colors: 40, 40, 40, 40
			        5235 => x"00000000",		-- colors: 40, 40, 40, 40
			        5236 => x"00000000",		-- colors: 40, 40, 40, 40
			        5237 => x"00000000",		-- colors: 40, 40, 40, 40
			        5238 => x"00000000",		-- colors: 40, 40, 40, 40
			        5239 => x"00000000",		-- colors: 40, 40, 40, 40
			        5240 => x"00000000",		-- colors: 40, 40, 40, 40
			        5241 => x"00000000",		-- colors: 40, 40, 40, 40
			        5242 => x"00000000",		-- colors: 40, 40, 40, 40
			        5243 => x"00000000",		-- colors: 40, 40, 40, 40
			        5244 => x"00000000",		-- colors: 40, 40, 40, 40
			        5245 => x"00000000",		-- colors: 40, 40, 40, 40
			        5246 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 78
			        5247 => x"00000000",		-- colors: 40, 40, 40, 40
			        5248 => x"00000000",		-- colors: 40, 40, 40, 40
			        5249 => x"00000000",		-- colors: 40, 40, 40, 40
			        5250 => x"00000000",		-- colors: 40, 40, 40, 40
			        5251 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5252 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5253 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5254 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5255 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5256 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5257 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5258 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5259 => x"00000000",		-- colors: 40, 40, 40, 40
			        5260 => x"00000000",		-- colors: 40, 40, 40, 40
			        5261 => x"00000000",		-- colors: 40, 40, 40, 40
			        5262 => x"00000000",		-- colors: 40, 40, 40, 40
			        5263 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5264 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5265 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5266 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5267 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5268 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5269 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5270 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5271 => x"00000000",		-- colors: 40, 40, 40, 40
			        5272 => x"00000000",		-- colors: 40, 40, 40, 40
			        5273 => x"00000000",		-- colors: 40, 40, 40, 40
			        5274 => x"00000000",		-- colors: 40, 40, 40, 40
			        5275 => x"00000000",		-- colors: 40, 40, 40, 40
			        5276 => x"00000000",		-- colors: 40, 40, 40, 40
			        5277 => x"00000000",		-- colors: 40, 40, 40, 40
			        5278 => x"00000000",		-- colors: 40, 40, 40, 40
			        5279 => x"00000000",		-- colors: 40, 40, 40, 40
			        5280 => x"00000000",		-- colors: 40, 40, 40, 40
			        5281 => x"00000000",		-- colors: 40, 40, 40, 40
			        5282 => x"00000000",		-- colors: 40, 40, 40, 40
			        5283 => x"00000000",		-- colors: 40, 40, 40, 40
			        5284 => x"00000000",		-- colors: 40, 40, 40, 40
			        5285 => x"00000000",		-- colors: 40, 40, 40, 40
			        5286 => x"00000000",		-- colors: 40, 40, 40, 40
			        5287 => x"00000000",		-- colors: 40, 40, 40, 40
			        5288 => x"00000000",		-- colors: 40, 40, 40, 40
			        5289 => x"00000000",		-- colors: 40, 40, 40, 40
			        5290 => x"00000000",		-- colors: 40, 40, 40, 40
			        5291 => x"00000000",		-- colors: 40, 40, 40, 40
			        5292 => x"00000000",		-- colors: 40, 40, 40, 40
			        5293 => x"00000000",		-- colors: 40, 40, 40, 40
			        5294 => x"00000000",		-- colors: 40, 40, 40, 40
			        5295 => x"00000000",		-- colors: 40, 40, 40, 40
			        5296 => x"00000000",		-- colors: 40, 40, 40, 40
			        5297 => x"00000000",		-- colors: 40, 40, 40, 40
			        5298 => x"00000000",		-- colors: 40, 40, 40, 40
			        5299 => x"00000000",		-- colors: 40, 40, 40, 40
			        5300 => x"00000000",		-- colors: 40, 40, 40, 40
			        5301 => x"00000000",		-- colors: 40, 40, 40, 40
			        5302 => x"00000000",		-- colors: 40, 40, 40, 40
			        5303 => x"00000000",		-- colors: 40, 40, 40, 40
			        5304 => x"00000000",		-- colors: 40, 40, 40, 40
			        5305 => x"00000000",		-- colors: 40, 40, 40, 40
			        5306 => x"00000000",		-- colors: 40, 40, 40, 40
			        5307 => x"00000000",		-- colors: 40, 40, 40, 40
			        5308 => x"00000000",		-- colors: 40, 40, 40, 40
			        5309 => x"00000000",		-- colors: 40, 40, 40, 40
			        5310 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 79
			        5311 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5312 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5313 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5314 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5315 => x"00000000",		-- colors: 40, 40, 40, 40
			        5316 => x"00000000",		-- colors: 40, 40, 40, 40
			        5317 => x"00000000",		-- colors: 40, 40, 40, 40
			        5318 => x"00000000",		-- colors: 40, 40, 40, 40
			        5319 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5320 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5321 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5322 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5323 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5324 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5325 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5326 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5327 => x"00000000",		-- colors: 40, 40, 40, 40
			        5328 => x"00000000",		-- colors: 40, 40, 40, 40
			        5329 => x"00000000",		-- colors: 40, 40, 40, 40
			        5330 => x"00000000",		-- colors: 40, 40, 40, 40
			        5331 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5332 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5333 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5334 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5335 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5336 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5337 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5338 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5339 => x"00000000",		-- colors: 40, 40, 40, 40
			        5340 => x"00000000",		-- colors: 40, 40, 40, 40
			        5341 => x"00000000",		-- colors: 40, 40, 40, 40
			        5342 => x"00000000",		-- colors: 40, 40, 40, 40
			        5343 => x"00000000",		-- colors: 40, 40, 40, 40
			        5344 => x"00000000",		-- colors: 40, 40, 40, 40
			        5345 => x"00000000",		-- colors: 40, 40, 40, 40
			        5346 => x"00000000",		-- colors: 40, 40, 40, 40
			        5347 => x"00000000",		-- colors: 40, 40, 40, 40
			        5348 => x"00000000",		-- colors: 40, 40, 40, 40
			        5349 => x"00000000",		-- colors: 40, 40, 40, 40
			        5350 => x"00000000",		-- colors: 40, 40, 40, 40
			        5351 => x"00000000",		-- colors: 40, 40, 40, 40
			        5352 => x"00000000",		-- colors: 40, 40, 40, 40
			        5353 => x"00000000",		-- colors: 40, 40, 40, 40
			        5354 => x"00000000",		-- colors: 40, 40, 40, 40
			        5355 => x"00000000",		-- colors: 40, 40, 40, 40
			        5356 => x"00000000",		-- colors: 40, 40, 40, 40
			        5357 => x"00000000",		-- colors: 40, 40, 40, 40
			        5358 => x"00000000",		-- colors: 40, 40, 40, 40
			        5359 => x"00000000",		-- colors: 40, 40, 40, 40
			        5360 => x"00000000",		-- colors: 40, 40, 40, 40
			        5361 => x"00000000",		-- colors: 40, 40, 40, 40
			        5362 => x"00000000",		-- colors: 40, 40, 40, 40
			        5363 => x"00000000",		-- colors: 40, 40, 40, 40
			        5364 => x"00000000",		-- colors: 40, 40, 40, 40
			        5365 => x"00000000",		-- colors: 40, 40, 40, 40
			        5366 => x"00000000",		-- colors: 40, 40, 40, 40
			        5367 => x"00000000",		-- colors: 40, 40, 40, 40
			        5368 => x"00000000",		-- colors: 40, 40, 40, 40
			        5369 => x"00000000",		-- colors: 40, 40, 40, 40
			        5370 => x"00000000",		-- colors: 40, 40, 40, 40
			        5371 => x"00000000",		-- colors: 40, 40, 40, 40
			        5372 => x"00000000",		-- colors: 40, 40, 40, 40
			        5373 => x"00000000",		-- colors: 40, 40, 40, 40
			        5374 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 80
			        5375 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5376 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5377 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5378 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5379 => x"00000000",		-- colors: 40, 40, 40, 40
			        5380 => x"00000000",		-- colors: 40, 40, 40, 40
			        5381 => x"00000000",		-- colors: 40, 40, 40, 40
			        5382 => x"00000000",		-- colors: 40, 40, 40, 40
			        5383 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5384 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5385 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5386 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5387 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5388 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5389 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5390 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5391 => x"00000000",		-- colors: 40, 40, 40, 40
			        5392 => x"00000000",		-- colors: 40, 40, 40, 40
			        5393 => x"00000000",		-- colors: 40, 40, 40, 40
			        5394 => x"00000000",		-- colors: 40, 40, 40, 40
			        5395 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5396 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5397 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5398 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5399 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5400 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5401 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5402 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5403 => x"00000000",		-- colors: 40, 40, 40, 40
			        5404 => x"00000000",		-- colors: 40, 40, 40, 40
			        5405 => x"00000000",		-- colors: 40, 40, 40, 40
			        5406 => x"00000000",		-- colors: 40, 40, 40, 40
			        5407 => x"00000000",		-- colors: 40, 40, 40, 40
			        5408 => x"00000000",		-- colors: 40, 40, 40, 40
			        5409 => x"00000000",		-- colors: 40, 40, 40, 40
			        5410 => x"00000000",		-- colors: 40, 40, 40, 40
			        5411 => x"00000000",		-- colors: 40, 40, 40, 40
			        5412 => x"00000000",		-- colors: 40, 40, 40, 40
			        5413 => x"00000000",		-- colors: 40, 40, 40, 40
			        5414 => x"00000000",		-- colors: 40, 40, 40, 40
			        5415 => x"00000000",		-- colors: 40, 40, 40, 40
			        5416 => x"00000000",		-- colors: 40, 40, 40, 40
			        5417 => x"00000000",		-- colors: 40, 40, 40, 40
			        5418 => x"00000000",		-- colors: 40, 40, 40, 40
			        5419 => x"00000000",		-- colors: 40, 40, 40, 40
			        5420 => x"00000000",		-- colors: 40, 40, 40, 40
			        5421 => x"00000000",		-- colors: 40, 40, 40, 40
			        5422 => x"00000000",		-- colors: 40, 40, 40, 40
			        5423 => x"00000000",		-- colors: 40, 40, 40, 40
			        5424 => x"00000000",		-- colors: 40, 40, 40, 40
			        5425 => x"00000000",		-- colors: 40, 40, 40, 40
			        5426 => x"00000000",		-- colors: 40, 40, 40, 40
			        5427 => x"00000000",		-- colors: 40, 40, 40, 40
			        5428 => x"00000000",		-- colors: 40, 40, 40, 40
			        5429 => x"00000000",		-- colors: 40, 40, 40, 40
			        5430 => x"00000000",		-- colors: 40, 40, 40, 40
			        5431 => x"00000000",		-- colors: 40, 40, 40, 40
			        5432 => x"00000000",		-- colors: 40, 40, 40, 40
			        5433 => x"00000000",		-- colors: 40, 40, 40, 40
			        5434 => x"00000000",		-- colors: 40, 40, 40, 40
			        5435 => x"00000000",		-- colors: 40, 40, 40, 40
			        5436 => x"00000000",		-- colors: 40, 40, 40, 40
			        5437 => x"00000000",		-- colors: 40, 40, 40, 40
			        5438 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 81
			        5439 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5440 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5441 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5442 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5443 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5444 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5445 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5446 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5447 => x"00000000",		-- colors: 40, 40, 40, 40
			        5448 => x"00000000",		-- colors: 40, 40, 40, 40
			        5449 => x"00000000",		-- colors: 40, 40, 40, 40
			        5450 => x"00000000",		-- colors: 40, 40, 40, 40
			        5451 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5452 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5453 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5454 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5455 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5456 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5457 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5458 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5459 => x"00000000",		-- colors: 40, 40, 40, 40
			        5460 => x"00000000",		-- colors: 40, 40, 40, 40
			        5461 => x"00000000",		-- colors: 40, 40, 40, 40
			        5462 => x"00000000",		-- colors: 40, 40, 40, 40
			        5463 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5464 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5465 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5466 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5467 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5468 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5469 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5470 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5471 => x"00000000",		-- colors: 40, 40, 40, 40
			        5472 => x"00000000",		-- colors: 40, 40, 40, 40
			        5473 => x"00000000",		-- colors: 40, 40, 40, 40
			        5474 => x"00000000",		-- colors: 40, 40, 40, 40
			        5475 => x"00000000",		-- colors: 40, 40, 40, 40
			        5476 => x"00000000",		-- colors: 40, 40, 40, 40
			        5477 => x"00000000",		-- colors: 40, 40, 40, 40
			        5478 => x"00000000",		-- colors: 40, 40, 40, 40
			        5479 => x"00000000",		-- colors: 40, 40, 40, 40
			        5480 => x"00000000",		-- colors: 40, 40, 40, 40
			        5481 => x"00000000",		-- colors: 40, 40, 40, 40
			        5482 => x"00000000",		-- colors: 40, 40, 40, 40
			        5483 => x"00000000",		-- colors: 40, 40, 40, 40
			        5484 => x"00000000",		-- colors: 40, 40, 40, 40
			        5485 => x"00000000",		-- colors: 40, 40, 40, 40
			        5486 => x"00000000",		-- colors: 40, 40, 40, 40
			        5487 => x"00000000",		-- colors: 40, 40, 40, 40
			        5488 => x"00000000",		-- colors: 40, 40, 40, 40
			        5489 => x"00000000",		-- colors: 40, 40, 40, 40
			        5490 => x"00000000",		-- colors: 40, 40, 40, 40
			        5491 => x"00000000",		-- colors: 40, 40, 40, 40
			        5492 => x"00000000",		-- colors: 40, 40, 40, 40
			        5493 => x"00000000",		-- colors: 40, 40, 40, 40
			        5494 => x"00000000",		-- colors: 40, 40, 40, 40
			        5495 => x"00000000",		-- colors: 40, 40, 40, 40
			        5496 => x"00000000",		-- colors: 40, 40, 40, 40
			        5497 => x"00000000",		-- colors: 40, 40, 40, 40
			        5498 => x"00000000",		-- colors: 40, 40, 40, 40
			        5499 => x"00000000",		-- colors: 40, 40, 40, 40
			        5500 => x"00000000",		-- colors: 40, 40, 40, 40
			        5501 => x"00000000",		-- colors: 40, 40, 40, 40
			        5502 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 82
			        5503 => x"00000000",		-- colors: 40, 40, 40, 40
			        5504 => x"00000000",		-- colors: 40, 40, 40, 40
			        5505 => x"00000000",		-- colors: 40, 40, 40, 40
			        5506 => x"00000000",		-- colors: 40, 40, 40, 40
			        5507 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5508 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5509 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5510 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5511 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5512 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5513 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5514 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5515 => x"00000000",		-- colors: 40, 40, 40, 40
			        5516 => x"00000000",		-- colors: 40, 40, 40, 40
			        5517 => x"00000000",		-- colors: 40, 40, 40, 40
			        5518 => x"00000000",		-- colors: 40, 40, 40, 40
			        5519 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5520 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5521 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5522 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5523 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5524 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5525 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5526 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5527 => x"00000000",		-- colors: 40, 40, 40, 40
			        5528 => x"00000000",		-- colors: 40, 40, 40, 40
			        5529 => x"00000000",		-- colors: 40, 40, 40, 40
			        5530 => x"00000000",		-- colors: 40, 40, 40, 40
			        5531 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5532 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5533 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5534 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5535 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5536 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5537 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5538 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5539 => x"00000000",		-- colors: 40, 40, 40, 40
			        5540 => x"00000000",		-- colors: 40, 40, 40, 40
			        5541 => x"00000000",		-- colors: 40, 40, 40, 40
			        5542 => x"00000000",		-- colors: 40, 40, 40, 40
			        5543 => x"32323232",		-- colors: 50, 50, 50, 50
			        5544 => x"32323232",		-- colors: 50, 50, 50, 50
			        5545 => x"32323232",		-- colors: 50, 50, 50, 50
			        5546 => x"32323232",		-- colors: 50, 50, 50, 50
			        5547 => x"00000000",		-- colors: 40, 40, 40, 40
			        5548 => x"00000000",		-- colors: 40, 40, 40, 40
			        5549 => x"00000000",		-- colors: 40, 40, 40, 40
			        5550 => x"00000000",		-- colors: 40, 40, 40, 40
			        5551 => x"00000000",		-- colors: 40, 40, 40, 40
			        5552 => x"00000000",		-- colors: 40, 40, 40, 40
			        5553 => x"00000000",		-- colors: 40, 40, 40, 40
			        5554 => x"00000000",		-- colors: 40, 40, 40, 40
			        5555 => x"00000000",		-- colors: 40, 40, 40, 40
			        5556 => x"00000000",		-- colors: 40, 40, 40, 40
			        5557 => x"00000000",		-- colors: 40, 40, 40, 40
			        5558 => x"00000000",		-- colors: 40, 40, 40, 40
			        5559 => x"32323232",		-- colors: 50, 50, 50, 50
			        5560 => x"32323232",		-- colors: 50, 50, 50, 50
			        5561 => x"32323232",		-- colors: 50, 50, 50, 50
			        5562 => x"32323232",		-- colors: 50, 50, 50, 50
			        5563 => x"00000000",		-- colors: 40, 40, 40, 40
			        5564 => x"00000000",		-- colors: 40, 40, 40, 40
			        5565 => x"00000000",		-- colors: 40, 40, 40, 40
			        5566 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 83
			        5567 => x"00000000",		-- colors: 40, 40, 40, 40
			        5568 => x"00000000",		-- colors: 40, 40, 40, 40
			        5569 => x"00000000",		-- colors: 40, 40, 40, 40
			        5570 => x"00000000",		-- colors: 40, 40, 40, 40
			        5571 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5572 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5573 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5574 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5575 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5576 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5577 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5578 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5579 => x"00000000",		-- colors: 40, 40, 40, 40
			        5580 => x"00000000",		-- colors: 40, 40, 40, 40
			        5581 => x"00000000",		-- colors: 40, 40, 40, 40
			        5582 => x"00000000",		-- colors: 40, 40, 40, 40
			        5583 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5584 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5585 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5586 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5587 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5588 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5589 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5590 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5591 => x"00000000",		-- colors: 40, 40, 40, 40
			        5592 => x"00000000",		-- colors: 40, 40, 40, 40
			        5593 => x"00000000",		-- colors: 40, 40, 40, 40
			        5594 => x"00000000",		-- colors: 40, 40, 40, 40
			        5595 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5596 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5597 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5598 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5599 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5600 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5601 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5602 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5603 => x"00000000",		-- colors: 40, 40, 40, 40
			        5604 => x"00000000",		-- colors: 40, 40, 40, 40
			        5605 => x"00000000",		-- colors: 40, 40, 40, 40
			        5606 => x"00000000",		-- colors: 40, 40, 40, 40
			        5607 => x"00000000",		-- colors: 40, 40, 40, 40
			        5608 => x"00000000",		-- colors: 40, 40, 40, 40
			        5609 => x"00000000",		-- colors: 40, 40, 40, 40
			        5610 => x"00000000",		-- colors: 40, 40, 40, 40
			        5611 => x"00000000",		-- colors: 40, 40, 40, 40
			        5612 => x"00000000",		-- colors: 40, 40, 40, 40
			        5613 => x"00000000",		-- colors: 40, 40, 40, 40
			        5614 => x"00000000",		-- colors: 40, 40, 40, 40
			        5615 => x"00000000",		-- colors: 40, 40, 40, 40
			        5616 => x"00000000",		-- colors: 40, 40, 40, 40
			        5617 => x"00000000",		-- colors: 40, 40, 40, 40
			        5618 => x"00000000",		-- colors: 40, 40, 40, 40
			        5619 => x"00000000",		-- colors: 40, 40, 40, 40
			        5620 => x"00000000",		-- colors: 40, 40, 40, 40
			        5621 => x"00000000",		-- colors: 40, 40, 40, 40
			        5622 => x"00000000",		-- colors: 40, 40, 40, 40
			        5623 => x"00000000",		-- colors: 40, 40, 40, 40
			        5624 => x"00000000",		-- colors: 40, 40, 40, 40
			        5625 => x"00000000",		-- colors: 40, 40, 40, 40
			        5626 => x"00000000",		-- colors: 40, 40, 40, 40
			        5627 => x"00000000",		-- colors: 40, 40, 40, 40
			        5628 => x"00000000",		-- colors: 40, 40, 40, 40
			        5629 => x"00000000",		-- colors: 40, 40, 40, 40
			        5630 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 84
			        5631 => x"00000000",		-- colors: 40, 40, 40, 40
			        5632 => x"00000000",		-- colors: 40, 40, 40, 40
			        5633 => x"00000000",		-- colors: 40, 40, 40, 40
			        5634 => x"00000000",		-- colors: 40, 40, 40, 40
			        5635 => x"00000000",		-- colors: 40, 40, 40, 40
			        5636 => x"00000000",		-- colors: 40, 40, 40, 40
			        5637 => x"00000000",		-- colors: 40, 40, 40, 40
			        5638 => x"00000000",		-- colors: 40, 40, 40, 40
			        5639 => x"00000000",		-- colors: 40, 40, 40, 40
			        5640 => x"00000000",		-- colors: 40, 40, 40, 40
			        5641 => x"00000000",		-- colors: 40, 40, 40, 40
			        5642 => x"00000000",		-- colors: 40, 40, 40, 40
			        5643 => x"00000000",		-- colors: 40, 40, 40, 40
			        5644 => x"00000000",		-- colors: 40, 40, 40, 40
			        5645 => x"00000000",		-- colors: 40, 40, 40, 40
			        5646 => x"00000000",		-- colors: 40, 40, 40, 40
			        5647 => x"00000000",		-- colors: 40, 40, 40, 40
			        5648 => x"00000000",		-- colors: 40, 40, 40, 40
			        5649 => x"00000000",		-- colors: 40, 40, 40, 40
			        5650 => x"00000000",		-- colors: 40, 40, 40, 40
			        5651 => x"00000000",		-- colors: 40, 40, 40, 40
			        5652 => x"00000000",		-- colors: 40, 40, 40, 40
			        5653 => x"00000000",		-- colors: 40, 40, 40, 40
			        5654 => x"00000000",		-- colors: 40, 40, 40, 40
			        5655 => x"00000000",		-- colors: 40, 40, 40, 40
			        5656 => x"00000000",		-- colors: 40, 40, 40, 40
			        5657 => x"00000000",		-- colors: 40, 40, 40, 40
			        5658 => x"00000000",		-- colors: 40, 40, 40, 40
			        5659 => x"00000000",		-- colors: 40, 40, 40, 40
			        5660 => x"00000000",		-- colors: 40, 40, 40, 40
			        5661 => x"00000000",		-- colors: 40, 40, 40, 40
			        5662 => x"00000000",		-- colors: 40, 40, 40, 40
			        5663 => x"00000000",		-- colors: 40, 40, 40, 40
			        5664 => x"00000000",		-- colors: 40, 40, 40, 40
			        5665 => x"00000000",		-- colors: 40, 40, 40, 40
			        5666 => x"00000000",		-- colors: 40, 40, 40, 40
			        5667 => x"00000000",		-- colors: 40, 40, 40, 40
			        5668 => x"00000000",		-- colors: 40, 40, 40, 40
			        5669 => x"00000000",		-- colors: 40, 40, 40, 40
			        5670 => x"00000000",		-- colors: 40, 40, 40, 40
			        5671 => x"00000000",		-- colors: 40, 40, 40, 40
			        5672 => x"00000000",		-- colors: 40, 40, 40, 40
			        5673 => x"00000000",		-- colors: 40, 40, 40, 40
			        5674 => x"00000000",		-- colors: 40, 40, 40, 40
			        5675 => x"00000000",		-- colors: 40, 40, 40, 40
			        5676 => x"00000000",		-- colors: 40, 40, 40, 40
			        5677 => x"00000000",		-- colors: 40, 40, 40, 40
			        5678 => x"00000000",		-- colors: 40, 40, 40, 40
			        5679 => x"00000000",		-- colors: 40, 40, 40, 40
			        5680 => x"00000000",		-- colors: 40, 40, 40, 40
			        5681 => x"00000000",		-- colors: 40, 40, 40, 40
			        5682 => x"00000000",		-- colors: 40, 40, 40, 40
			        5683 => x"00000000",		-- colors: 40, 40, 40, 40
			        5684 => x"00000000",		-- colors: 40, 40, 40, 40
			        5685 => x"00000000",		-- colors: 40, 40, 40, 40
			        5686 => x"00000000",		-- colors: 40, 40, 40, 40
			        5687 => x"00000000",		-- colors: 40, 40, 40, 40
			        5688 => x"00000000",		-- colors: 40, 40, 40, 40
			        5689 => x"00000000",		-- colors: 40, 40, 40, 40
			        5690 => x"00000000",		-- colors: 40, 40, 40, 40
			        5691 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5692 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5693 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5694 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60

			                --  sprite 85
			        5695 => x"00000000",		-- colors: 40, 40, 40, 40
			        5696 => x"00000000",		-- colors: 40, 40, 40, 40
			        5697 => x"00000000",		-- colors: 40, 40, 40, 40
			        5698 => x"00000000",		-- colors: 40, 40, 40, 40
			        5699 => x"00000000",		-- colors: 40, 40, 40, 40
			        5700 => x"00000000",		-- colors: 40, 40, 40, 40
			        5701 => x"00000000",		-- colors: 40, 40, 40, 40
			        5702 => x"00000000",		-- colors: 40, 40, 40, 40
			        5703 => x"00000000",		-- colors: 40, 40, 40, 40
			        5704 => x"00000000",		-- colors: 40, 40, 40, 40
			        5705 => x"00000000",		-- colors: 40, 40, 40, 40
			        5706 => x"00000000",		-- colors: 40, 40, 40, 40
			        5707 => x"00000000",		-- colors: 40, 40, 40, 40
			        5708 => x"00000000",		-- colors: 40, 40, 40, 40
			        5709 => x"00000000",		-- colors: 40, 40, 40, 40
			        5710 => x"00000000",		-- colors: 40, 40, 40, 40
			        5711 => x"00000000",		-- colors: 40, 40, 40, 40
			        5712 => x"00000000",		-- colors: 40, 40, 40, 40
			        5713 => x"00000000",		-- colors: 40, 40, 40, 40
			        5714 => x"00000000",		-- colors: 40, 40, 40, 40
			        5715 => x"00000000",		-- colors: 40, 40, 40, 40
			        5716 => x"00000000",		-- colors: 40, 40, 40, 40
			        5717 => x"00000000",		-- colors: 40, 40, 40, 40
			        5718 => x"00000000",		-- colors: 40, 40, 40, 40
			        5719 => x"00000000",		-- colors: 40, 40, 40, 40
			        5720 => x"00000000",		-- colors: 40, 40, 40, 40
			        5721 => x"00000000",		-- colors: 40, 40, 40, 40
			        5722 => x"00000000",		-- colors: 40, 40, 40, 40
			        5723 => x"00000000",		-- colors: 40, 40, 40, 40
			        5724 => x"00000000",		-- colors: 40, 40, 40, 40
			        5725 => x"00000000",		-- colors: 40, 40, 40, 40
			        5726 => x"00000000",		-- colors: 40, 40, 40, 40
			        5727 => x"00000000",		-- colors: 40, 40, 40, 40
			        5728 => x"00000000",		-- colors: 40, 40, 40, 40
			        5729 => x"00000000",		-- colors: 40, 40, 40, 40
			        5730 => x"00000000",		-- colors: 40, 40, 40, 40
			        5731 => x"00000000",		-- colors: 40, 40, 40, 40
			        5732 => x"00000000",		-- colors: 40, 40, 40, 40
			        5733 => x"00000000",		-- colors: 40, 40, 40, 40
			        5734 => x"00000000",		-- colors: 40, 40, 40, 40
			        5735 => x"00000000",		-- colors: 40, 40, 40, 40
			        5736 => x"00000000",		-- colors: 40, 40, 40, 40
			        5737 => x"00000000",		-- colors: 40, 40, 40, 40
			        5738 => x"00000000",		-- colors: 40, 40, 40, 40
			        5739 => x"00000000",		-- colors: 40, 40, 40, 40
			        5740 => x"00000000",		-- colors: 40, 40, 40, 40
			        5741 => x"00000000",		-- colors: 40, 40, 40, 40
			        5742 => x"00000000",		-- colors: 40, 40, 40, 40
			        5743 => x"00000000",		-- colors: 40, 40, 40, 40
			        5744 => x"00000000",		-- colors: 40, 40, 40, 40
			        5745 => x"00000000",		-- colors: 40, 40, 40, 40
			        5746 => x"00000000",		-- colors: 40, 40, 40, 40
			        5747 => x"00000000",		-- colors: 40, 40, 40, 40
			        5748 => x"00000000",		-- colors: 40, 40, 40, 40
			        5749 => x"00000000",		-- colors: 40, 40, 40, 40
			        5750 => x"00000000",		-- colors: 40, 40, 40, 40
			        5751 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5752 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5753 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5754 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5755 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5756 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5757 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5758 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60

			                --  sprite 86
			        5759 => x"00000000",		-- colors: 40, 40, 40, 40
			        5760 => x"00000000",		-- colors: 40, 40, 40, 40
			        5761 => x"00000000",		-- colors: 40, 40, 40, 40
			        5762 => x"00000000",		-- colors: 40, 40, 40, 40
			        5763 => x"00000000",		-- colors: 40, 40, 40, 40
			        5764 => x"00000000",		-- colors: 40, 40, 40, 40
			        5765 => x"00000000",		-- colors: 40, 40, 40, 40
			        5766 => x"00000000",		-- colors: 40, 40, 40, 40
			        5767 => x"00000000",		-- colors: 40, 40, 40, 40
			        5768 => x"00000000",		-- colors: 40, 40, 40, 40
			        5769 => x"00000000",		-- colors: 40, 40, 40, 40
			        5770 => x"00000000",		-- colors: 40, 40, 40, 40
			        5771 => x"00000000",		-- colors: 40, 40, 40, 40
			        5772 => x"00000000",		-- colors: 40, 40, 40, 40
			        5773 => x"00000000",		-- colors: 40, 40, 40, 40
			        5774 => x"00000000",		-- colors: 40, 40, 40, 40
			        5775 => x"00000000",		-- colors: 40, 40, 40, 40
			        5776 => x"00000000",		-- colors: 40, 40, 40, 40
			        5777 => x"00000000",		-- colors: 40, 40, 40, 40
			        5778 => x"00000000",		-- colors: 40, 40, 40, 40
			        5779 => x"00000000",		-- colors: 40, 40, 40, 40
			        5780 => x"00000000",		-- colors: 40, 40, 40, 40
			        5781 => x"00000000",		-- colors: 40, 40, 40, 40
			        5782 => x"00000000",		-- colors: 40, 40, 40, 40
			        5783 => x"00000000",		-- colors: 40, 40, 40, 40
			        5784 => x"00000000",		-- colors: 40, 40, 40, 40
			        5785 => x"00000000",		-- colors: 40, 40, 40, 40
			        5786 => x"00000000",		-- colors: 40, 40, 40, 40
			        5787 => x"00000000",		-- colors: 40, 40, 40, 40
			        5788 => x"00000000",		-- colors: 40, 40, 40, 40
			        5789 => x"00000000",		-- colors: 40, 40, 40, 40
			        5790 => x"00000000",		-- colors: 40, 40, 40, 40
			        5791 => x"00000000",		-- colors: 40, 40, 40, 40
			        5792 => x"00000000",		-- colors: 40, 40, 40, 40
			        5793 => x"00000000",		-- colors: 40, 40, 40, 40
			        5794 => x"00000000",		-- colors: 40, 40, 40, 40
			        5795 => x"00000000",		-- colors: 40, 40, 40, 40
			        5796 => x"00000000",		-- colors: 40, 40, 40, 40
			        5797 => x"00000000",		-- colors: 40, 40, 40, 40
			        5798 => x"00000000",		-- colors: 40, 40, 40, 40
			        5799 => x"00000000",		-- colors: 40, 40, 40, 40
			        5800 => x"00000000",		-- colors: 40, 40, 40, 40
			        5801 => x"00000000",		-- colors: 40, 40, 40, 40
			        5802 => x"00000000",		-- colors: 40, 40, 40, 40
			        5803 => x"00000000",		-- colors: 40, 40, 40, 40
			        5804 => x"00000000",		-- colors: 40, 40, 40, 40
			        5805 => x"00000000",		-- colors: 40, 40, 40, 40
			        5806 => x"00000000",		-- colors: 40, 40, 40, 40
			        5807 => x"00000000",		-- colors: 40, 40, 40, 40
			        5808 => x"00000000",		-- colors: 40, 40, 40, 40
			        5809 => x"00000000",		-- colors: 40, 40, 40, 40
			        5810 => x"00000000",		-- colors: 40, 40, 40, 40
			        5811 => x"00000000",		-- colors: 40, 40, 40, 40
			        5812 => x"00000000",		-- colors: 40, 40, 40, 40
			        5813 => x"00000000",		-- colors: 40, 40, 40, 40
			        5814 => x"00000000",		-- colors: 40, 40, 40, 40
			        5815 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5816 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5817 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5818 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5819 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5820 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5821 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5822 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60

			                --  sprite 87
			        5823 => x"00000000",		-- colors: 40, 40, 40, 40
			        5824 => x"00000000",		-- colors: 40, 40, 40, 40
			        5825 => x"00000000",		-- colors: 40, 40, 40, 40
			        5826 => x"00000000",		-- colors: 40, 40, 40, 40
			        5827 => x"00000000",		-- colors: 40, 40, 40, 40
			        5828 => x"00000000",		-- colors: 40, 40, 40, 40
			        5829 => x"00000000",		-- colors: 40, 40, 40, 40
			        5830 => x"00000000",		-- colors: 40, 40, 40, 40
			        5831 => x"00000000",		-- colors: 40, 40, 40, 40
			        5832 => x"00000000",		-- colors: 40, 40, 40, 40
			        5833 => x"00000000",		-- colors: 40, 40, 40, 40
			        5834 => x"00000000",		-- colors: 40, 40, 40, 40
			        5835 => x"00000000",		-- colors: 40, 40, 40, 40
			        5836 => x"00000000",		-- colors: 40, 40, 40, 40
			        5837 => x"00000000",		-- colors: 40, 40, 40, 40
			        5838 => x"00000000",		-- colors: 40, 40, 40, 40
			        5839 => x"00000000",		-- colors: 40, 40, 40, 40
			        5840 => x"00000000",		-- colors: 40, 40, 40, 40
			        5841 => x"00000000",		-- colors: 40, 40, 40, 40
			        5842 => x"00000000",		-- colors: 40, 40, 40, 40
			        5843 => x"00000000",		-- colors: 40, 40, 40, 40
			        5844 => x"00000000",		-- colors: 40, 40, 40, 40
			        5845 => x"00000000",		-- colors: 40, 40, 40, 40
			        5846 => x"00000000",		-- colors: 40, 40, 40, 40
			        5847 => x"00000000",		-- colors: 40, 40, 40, 40
			        5848 => x"00000000",		-- colors: 40, 40, 40, 40
			        5849 => x"00000000",		-- colors: 40, 40, 40, 40
			        5850 => x"00000000",		-- colors: 40, 40, 40, 40
			        5851 => x"00000000",		-- colors: 40, 40, 40, 40
			        5852 => x"00000000",		-- colors: 40, 40, 40, 40
			        5853 => x"00000000",		-- colors: 40, 40, 40, 40
			        5854 => x"00000000",		-- colors: 40, 40, 40, 40
			        5855 => x"00000000",		-- colors: 40, 40, 40, 40
			        5856 => x"00000000",		-- colors: 40, 40, 40, 40
			        5857 => x"00000000",		-- colors: 40, 40, 40, 40
			        5858 => x"00000000",		-- colors: 40, 40, 40, 40
			        5859 => x"00000000",		-- colors: 40, 40, 40, 40
			        5860 => x"00000000",		-- colors: 40, 40, 40, 40
			        5861 => x"00000000",		-- colors: 40, 40, 40, 40
			        5862 => x"00000000",		-- colors: 40, 40, 40, 40
			        5863 => x"00000000",		-- colors: 40, 40, 40, 40
			        5864 => x"00000000",		-- colors: 40, 40, 40, 40
			        5865 => x"00000000",		-- colors: 40, 40, 40, 40
			        5866 => x"00000000",		-- colors: 40, 40, 40, 40
			        5867 => x"00000000",		-- colors: 40, 40, 40, 40
			        5868 => x"00000000",		-- colors: 40, 40, 40, 40
			        5869 => x"00000000",		-- colors: 40, 40, 40, 40
			        5870 => x"00000000",		-- colors: 40, 40, 40, 40
			        5871 => x"00000000",		-- colors: 40, 40, 40, 40
			        5872 => x"00000000",		-- colors: 40, 40, 40, 40
			        5873 => x"00000000",		-- colors: 40, 40, 40, 40
			        5874 => x"00000000",		-- colors: 40, 40, 40, 40
			        5875 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5876 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5877 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5878 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5879 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5880 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5881 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5882 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5883 => x"00000000",		-- colors: 40, 40, 40, 40
			        5884 => x"00000000",		-- colors: 40, 40, 40, 40
			        5885 => x"00000000",		-- colors: 40, 40, 40, 40
			        5886 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 88
			        5887 => x"00000000",		-- colors: 40, 40, 40, 40
			        5888 => x"00000000",		-- colors: 40, 40, 40, 40
			        5889 => x"00000000",		-- colors: 40, 40, 40, 40
			        5890 => x"00000000",		-- colors: 40, 40, 40, 40
			        5891 => x"00000000",		-- colors: 40, 40, 40, 40
			        5892 => x"00000000",		-- colors: 40, 40, 40, 40
			        5893 => x"00000000",		-- colors: 40, 40, 40, 40
			        5894 => x"00000000",		-- colors: 40, 40, 40, 40
			        5895 => x"00000000",		-- colors: 40, 40, 40, 40
			        5896 => x"00000000",		-- colors: 40, 40, 40, 40
			        5897 => x"00000000",		-- colors: 40, 40, 40, 40
			        5898 => x"00000000",		-- colors: 40, 40, 40, 40
			        5899 => x"00000000",		-- colors: 40, 40, 40, 40
			        5900 => x"00000000",		-- colors: 40, 40, 40, 40
			        5901 => x"00000000",		-- colors: 40, 40, 40, 40
			        5902 => x"00000000",		-- colors: 40, 40, 40, 40
			        5903 => x"00000000",		-- colors: 40, 40, 40, 40
			        5904 => x"00000000",		-- colors: 40, 40, 40, 40
			        5905 => x"00000000",		-- colors: 40, 40, 40, 40
			        5906 => x"00000000",		-- colors: 40, 40, 40, 40
			        5907 => x"00000000",		-- colors: 40, 40, 40, 40
			        5908 => x"00000000",		-- colors: 40, 40, 40, 40
			        5909 => x"00000000",		-- colors: 40, 40, 40, 40
			        5910 => x"00000000",		-- colors: 40, 40, 40, 40
			        5911 => x"00000000",		-- colors: 40, 40, 40, 40
			        5912 => x"00000000",		-- colors: 40, 40, 40, 40
			        5913 => x"00000000",		-- colors: 40, 40, 40, 40
			        5914 => x"00000000",		-- colors: 40, 40, 40, 40
			        5915 => x"00000000",		-- colors: 40, 40, 40, 40
			        5916 => x"00000000",		-- colors: 40, 40, 40, 40
			        5917 => x"00000000",		-- colors: 40, 40, 40, 40
			        5918 => x"00000000",		-- colors: 40, 40, 40, 40
			        5919 => x"00000000",		-- colors: 40, 40, 40, 40
			        5920 => x"00000000",		-- colors: 40, 40, 40, 40
			        5921 => x"00000000",		-- colors: 40, 40, 40, 40
			        5922 => x"00000000",		-- colors: 40, 40, 40, 40
			        5923 => x"00000000",		-- colors: 40, 40, 40, 40
			        5924 => x"00000000",		-- colors: 40, 40, 40, 40
			        5925 => x"00000000",		-- colors: 40, 40, 40, 40
			        5926 => x"00000000",		-- colors: 40, 40, 40, 40
			        5927 => x"00000000",		-- colors: 40, 40, 40, 40
			        5928 => x"00000000",		-- colors: 40, 40, 40, 40
			        5929 => x"00000000",		-- colors: 40, 40, 40, 40
			        5930 => x"00000000",		-- colors: 40, 40, 40, 40
			        5931 => x"00000000",		-- colors: 40, 40, 40, 40
			        5932 => x"00000000",		-- colors: 40, 40, 40, 40
			        5933 => x"00000000",		-- colors: 40, 40, 40, 40
			        5934 => x"00000000",		-- colors: 40, 40, 40, 40
			        5935 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5936 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5937 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5938 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5939 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5940 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5941 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5942 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5943 => x"00000000",		-- colors: 40, 40, 40, 40
			        5944 => x"00000000",		-- colors: 40, 40, 40, 40
			        5945 => x"00000000",		-- colors: 40, 40, 40, 40
			        5946 => x"00000000",		-- colors: 40, 40, 40, 40
			        5947 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5948 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5949 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        5950 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60

			                --  sprite 89
			        5951 => x"00000000",		-- colors: 40, 40, 40, 40
			        5952 => x"00000000",		-- colors: 40, 40, 40, 40
			        5953 => x"00000000",		-- colors: 40, 40, 40, 40
			        5954 => x"00000000",		-- colors: 40, 40, 40, 40
			        5955 => x"00000000",		-- colors: 40, 40, 40, 40
			        5956 => x"00000000",		-- colors: 40, 40, 40, 40
			        5957 => x"00000000",		-- colors: 40, 40, 40, 40
			        5958 => x"00000000",		-- colors: 40, 40, 40, 40
			        5959 => x"00000000",		-- colors: 40, 40, 40, 40
			        5960 => x"00000000",		-- colors: 40, 40, 40, 40
			        5961 => x"00000000",		-- colors: 40, 40, 40, 40
			        5962 => x"00000000",		-- colors: 40, 40, 40, 40
			        5963 => x"00000000",		-- colors: 40, 40, 40, 40
			        5964 => x"00000000",		-- colors: 40, 40, 40, 40
			        5965 => x"00000000",		-- colors: 40, 40, 40, 40
			        5966 => x"00000000",		-- colors: 40, 40, 40, 40
			        5967 => x"00000000",		-- colors: 40, 40, 40, 40
			        5968 => x"00000000",		-- colors: 40, 40, 40, 40
			        5969 => x"00000000",		-- colors: 40, 40, 40, 40
			        5970 => x"00000000",		-- colors: 40, 40, 40, 40
			        5971 => x"00000000",		-- colors: 40, 40, 40, 40
			        5972 => x"00000000",		-- colors: 40, 40, 40, 40
			        5973 => x"00000000",		-- colors: 40, 40, 40, 40
			        5974 => x"00000000",		-- colors: 40, 40, 40, 40
			        5975 => x"00000000",		-- colors: 40, 40, 40, 40
			        5976 => x"00000000",		-- colors: 40, 40, 40, 40
			        5977 => x"00000000",		-- colors: 40, 40, 40, 40
			        5978 => x"00000000",		-- colors: 40, 40, 40, 40
			        5979 => x"00000000",		-- colors: 40, 40, 40, 40
			        5980 => x"00000000",		-- colors: 40, 40, 40, 40
			        5981 => x"00000000",		-- colors: 40, 40, 40, 40
			        5982 => x"00000000",		-- colors: 40, 40, 40, 40
			        5983 => x"00000000",		-- colors: 40, 40, 40, 40
			        5984 => x"00000000",		-- colors: 40, 40, 40, 40
			        5985 => x"00000000",		-- colors: 40, 40, 40, 40
			        5986 => x"00000000",		-- colors: 40, 40, 40, 40
			        5987 => x"00000000",		-- colors: 40, 40, 40, 40
			        5988 => x"00000000",		-- colors: 40, 40, 40, 40
			        5989 => x"00000000",		-- colors: 40, 40, 40, 40
			        5990 => x"00000000",		-- colors: 40, 40, 40, 40
			        5991 => x"00000000",		-- colors: 40, 40, 40, 40
			        5992 => x"00000000",		-- colors: 40, 40, 40, 40
			        5993 => x"00000000",		-- colors: 40, 40, 40, 40
			        5994 => x"00000000",		-- colors: 40, 40, 40, 40
			        5995 => x"00000000",		-- colors: 40, 40, 40, 40
			        5996 => x"00000000",		-- colors: 40, 40, 40, 40
			        5997 => x"00000000",		-- colors: 40, 40, 40, 40
			        5998 => x"00000000",		-- colors: 40, 40, 40, 40
			        5999 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6000 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6001 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6002 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6003 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6004 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6005 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6006 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6007 => x"00000000",		-- colors: 40, 40, 40, 40
			        6008 => x"00000000",		-- colors: 40, 40, 40, 40
			        6009 => x"00000000",		-- colors: 40, 40, 40, 40
			        6010 => x"00000000",		-- colors: 40, 40, 40, 40
			        6011 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6012 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6013 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6014 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60

			                --  sprite 90
			        6015 => x"00000000",		-- colors: 40, 40, 40, 40
			        6016 => x"00000000",		-- colors: 40, 40, 40, 40
			        6017 => x"00000000",		-- colors: 40, 40, 40, 40
			        6018 => x"00000000",		-- colors: 40, 40, 40, 40
			        6019 => x"00000000",		-- colors: 40, 40, 40, 40
			        6020 => x"00000000",		-- colors: 40, 40, 40, 40
			        6021 => x"00000000",		-- colors: 40, 40, 40, 40
			        6022 => x"00000000",		-- colors: 40, 40, 40, 40
			        6023 => x"00000000",		-- colors: 40, 40, 40, 40
			        6024 => x"00000000",		-- colors: 40, 40, 40, 40
			        6025 => x"00000000",		-- colors: 40, 40, 40, 40
			        6026 => x"00000000",		-- colors: 40, 40, 40, 40
			        6027 => x"00000000",		-- colors: 40, 40, 40, 40
			        6028 => x"00000000",		-- colors: 40, 40, 40, 40
			        6029 => x"00000000",		-- colors: 40, 40, 40, 40
			        6030 => x"00000000",		-- colors: 40, 40, 40, 40
			        6031 => x"00000000",		-- colors: 40, 40, 40, 40
			        6032 => x"00000000",		-- colors: 40, 40, 40, 40
			        6033 => x"00000000",		-- colors: 40, 40, 40, 40
			        6034 => x"00000000",		-- colors: 40, 40, 40, 40
			        6035 => x"00000000",		-- colors: 40, 40, 40, 40
			        6036 => x"00000000",		-- colors: 40, 40, 40, 40
			        6037 => x"00000000",		-- colors: 40, 40, 40, 40
			        6038 => x"00000000",		-- colors: 40, 40, 40, 40
			        6039 => x"00000000",		-- colors: 40, 40, 40, 40
			        6040 => x"00000000",		-- colors: 40, 40, 40, 40
			        6041 => x"00000000",		-- colors: 40, 40, 40, 40
			        6042 => x"00000000",		-- colors: 40, 40, 40, 40
			        6043 => x"00000000",		-- colors: 40, 40, 40, 40
			        6044 => x"00000000",		-- colors: 40, 40, 40, 40
			        6045 => x"00000000",		-- colors: 40, 40, 40, 40
			        6046 => x"00000000",		-- colors: 40, 40, 40, 40
			        6047 => x"00000000",		-- colors: 40, 40, 40, 40
			        6048 => x"00000000",		-- colors: 40, 40, 40, 40
			        6049 => x"00000000",		-- colors: 40, 40, 40, 40
			        6050 => x"00000000",		-- colors: 40, 40, 40, 40
			        6051 => x"00000000",		-- colors: 40, 40, 40, 40
			        6052 => x"00000000",		-- colors: 40, 40, 40, 40
			        6053 => x"00000000",		-- colors: 40, 40, 40, 40
			        6054 => x"00000000",		-- colors: 40, 40, 40, 40
			        6055 => x"00000000",		-- colors: 40, 40, 40, 40
			        6056 => x"00000000",		-- colors: 40, 40, 40, 40
			        6057 => x"00000000",		-- colors: 40, 40, 40, 40
			        6058 => x"00000000",		-- colors: 40, 40, 40, 40
			        6059 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6060 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6061 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6062 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6063 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6064 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6065 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6066 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6067 => x"00000000",		-- colors: 40, 40, 40, 40
			        6068 => x"00000000",		-- colors: 40, 40, 40, 40
			        6069 => x"00000000",		-- colors: 40, 40, 40, 40
			        6070 => x"00000000",		-- colors: 40, 40, 40, 40
			        6071 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6072 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6073 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6074 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6075 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6076 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6077 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6078 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60

			                --  sprite 91
			        6079 => x"00000000",		-- colors: 40, 40, 40, 40
			        6080 => x"00000000",		-- colors: 40, 40, 40, 40
			        6081 => x"00000000",		-- colors: 40, 40, 40, 40
			        6082 => x"00000000",		-- colors: 40, 40, 40, 40
			        6083 => x"00000000",		-- colors: 40, 40, 40, 40
			        6084 => x"00000000",		-- colors: 40, 40, 40, 40
			        6085 => x"00000000",		-- colors: 40, 40, 40, 40
			        6086 => x"00000000",		-- colors: 40, 40, 40, 40
			        6087 => x"00000000",		-- colors: 40, 40, 40, 40
			        6088 => x"00000000",		-- colors: 40, 40, 40, 40
			        6089 => x"00000000",		-- colors: 40, 40, 40, 40
			        6090 => x"00000000",		-- colors: 40, 40, 40, 40
			        6091 => x"00000000",		-- colors: 40, 40, 40, 40
			        6092 => x"00000000",		-- colors: 40, 40, 40, 40
			        6093 => x"00000000",		-- colors: 40, 40, 40, 40
			        6094 => x"00000000",		-- colors: 40, 40, 40, 40
			        6095 => x"00000000",		-- colors: 40, 40, 40, 40
			        6096 => x"00000000",		-- colors: 40, 40, 40, 40
			        6097 => x"00000000",		-- colors: 40, 40, 40, 40
			        6098 => x"00000000",		-- colors: 40, 40, 40, 40
			        6099 => x"00000000",		-- colors: 40, 40, 40, 40
			        6100 => x"00000000",		-- colors: 40, 40, 40, 40
			        6101 => x"00000000",		-- colors: 40, 40, 40, 40
			        6102 => x"00000000",		-- colors: 40, 40, 40, 40
			        6103 => x"00000000",		-- colors: 40, 40, 40, 40
			        6104 => x"00000000",		-- colors: 40, 40, 40, 40
			        6105 => x"00000000",		-- colors: 40, 40, 40, 40
			        6106 => x"00000000",		-- colors: 40, 40, 40, 40
			        6107 => x"00000000",		-- colors: 40, 40, 40, 40
			        6108 => x"00000000",		-- colors: 40, 40, 40, 40
			        6109 => x"00000000",		-- colors: 40, 40, 40, 40
			        6110 => x"00000000",		-- colors: 40, 40, 40, 40
			        6111 => x"00000000",		-- colors: 40, 40, 40, 40
			        6112 => x"00000000",		-- colors: 40, 40, 40, 40
			        6113 => x"00000000",		-- colors: 40, 40, 40, 40
			        6114 => x"00000000",		-- colors: 40, 40, 40, 40
			        6115 => x"00000000",		-- colors: 40, 40, 40, 40
			        6116 => x"00000000",		-- colors: 40, 40, 40, 40
			        6117 => x"00000000",		-- colors: 40, 40, 40, 40
			        6118 => x"00000000",		-- colors: 40, 40, 40, 40
			        6119 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6120 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6121 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6122 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6123 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6124 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6125 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6126 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6127 => x"00000000",		-- colors: 40, 40, 40, 40
			        6128 => x"00000000",		-- colors: 40, 40, 40, 40
			        6129 => x"00000000",		-- colors: 40, 40, 40, 40
			        6130 => x"00000000",		-- colors: 40, 40, 40, 40
			        6131 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6132 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6133 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6134 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6135 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6136 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6137 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6138 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6139 => x"00000000",		-- colors: 40, 40, 40, 40
			        6140 => x"00000000",		-- colors: 40, 40, 40, 40
			        6141 => x"00000000",		-- colors: 40, 40, 40, 40
			        6142 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 92
			        6143 => x"00000000",		-- colors: 40, 40, 40, 40
			        6144 => x"00000000",		-- colors: 40, 40, 40, 40
			        6145 => x"00000000",		-- colors: 40, 40, 40, 40
			        6146 => x"00000000",		-- colors: 40, 40, 40, 40
			        6147 => x"00000000",		-- colors: 40, 40, 40, 40
			        6148 => x"00000000",		-- colors: 40, 40, 40, 40
			        6149 => x"00000000",		-- colors: 40, 40, 40, 40
			        6150 => x"00000000",		-- colors: 40, 40, 40, 40
			        6151 => x"00000000",		-- colors: 40, 40, 40, 40
			        6152 => x"00000000",		-- colors: 40, 40, 40, 40
			        6153 => x"00000000",		-- colors: 40, 40, 40, 40
			        6154 => x"00000000",		-- colors: 40, 40, 40, 40
			        6155 => x"00000000",		-- colors: 40, 40, 40, 40
			        6156 => x"00000000",		-- colors: 40, 40, 40, 40
			        6157 => x"00000000",		-- colors: 40, 40, 40, 40
			        6158 => x"00000000",		-- colors: 40, 40, 40, 40
			        6159 => x"00000000",		-- colors: 40, 40, 40, 40
			        6160 => x"00000000",		-- colors: 40, 40, 40, 40
			        6161 => x"00000000",		-- colors: 40, 40, 40, 40
			        6162 => x"00000000",		-- colors: 40, 40, 40, 40
			        6163 => x"00000000",		-- colors: 40, 40, 40, 40
			        6164 => x"00000000",		-- colors: 40, 40, 40, 40
			        6165 => x"00000000",		-- colors: 40, 40, 40, 40
			        6166 => x"00000000",		-- colors: 40, 40, 40, 40
			        6167 => x"00000000",		-- colors: 40, 40, 40, 40
			        6168 => x"00000000",		-- colors: 40, 40, 40, 40
			        6169 => x"00000000",		-- colors: 40, 40, 40, 40
			        6170 => x"00000000",		-- colors: 40, 40, 40, 40
			        6171 => x"00000000",		-- colors: 40, 40, 40, 40
			        6172 => x"00000000",		-- colors: 40, 40, 40, 40
			        6173 => x"00000000",		-- colors: 40, 40, 40, 40
			        6174 => x"00000000",		-- colors: 40, 40, 40, 40
			        6175 => x"00000000",		-- colors: 40, 40, 40, 40
			        6176 => x"00000000",		-- colors: 40, 40, 40, 40
			        6177 => x"00000000",		-- colors: 40, 40, 40, 40
			        6178 => x"00000000",		-- colors: 40, 40, 40, 40
			        6179 => x"00000000",		-- colors: 40, 40, 40, 40
			        6180 => x"00000000",		-- colors: 40, 40, 40, 40
			        6181 => x"00000000",		-- colors: 40, 40, 40, 40
			        6182 => x"00000000",		-- colors: 40, 40, 40, 40
			        6183 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6184 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6185 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6186 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6187 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6188 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6189 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6190 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6191 => x"00000000",		-- colors: 40, 40, 40, 40
			        6192 => x"00000000",		-- colors: 40, 40, 40, 40
			        6193 => x"00000000",		-- colors: 40, 40, 40, 40
			        6194 => x"00000000",		-- colors: 40, 40, 40, 40
			        6195 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6196 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6197 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6198 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6199 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6200 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6201 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6202 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6203 => x"00000000",		-- colors: 40, 40, 40, 40
			        6204 => x"00000000",		-- colors: 40, 40, 40, 40
			        6205 => x"00000000",		-- colors: 40, 40, 40, 40
			        6206 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 93
			        6207 => x"00000000",		-- colors: 40, 40, 40, 40
			        6208 => x"00000000",		-- colors: 40, 40, 40, 40
			        6209 => x"00000000",		-- colors: 40, 40, 40, 40
			        6210 => x"00000000",		-- colors: 40, 40, 40, 40
			        6211 => x"00000000",		-- colors: 40, 40, 40, 40
			        6212 => x"00000000",		-- colors: 40, 40, 40, 40
			        6213 => x"00000000",		-- colors: 40, 40, 40, 40
			        6214 => x"00000000",		-- colors: 40, 40, 40, 40
			        6215 => x"00000000",		-- colors: 40, 40, 40, 40
			        6216 => x"00000000",		-- colors: 40, 40, 40, 40
			        6217 => x"00000000",		-- colors: 40, 40, 40, 40
			        6218 => x"00000000",		-- colors: 40, 40, 40, 40
			        6219 => x"00000000",		-- colors: 40, 40, 40, 40
			        6220 => x"00000000",		-- colors: 40, 40, 40, 40
			        6221 => x"00000000",		-- colors: 40, 40, 40, 40
			        6222 => x"00000000",		-- colors: 40, 40, 40, 40
			        6223 => x"00000000",		-- colors: 40, 40, 40, 40
			        6224 => x"00000000",		-- colors: 40, 40, 40, 40
			        6225 => x"00000000",		-- colors: 40, 40, 40, 40
			        6226 => x"00000000",		-- colors: 40, 40, 40, 40
			        6227 => x"00000000",		-- colors: 40, 40, 40, 40
			        6228 => x"00000000",		-- colors: 40, 40, 40, 40
			        6229 => x"00000000",		-- colors: 40, 40, 40, 40
			        6230 => x"00000000",		-- colors: 40, 40, 40, 40
			        6231 => x"00000000",		-- colors: 40, 40, 40, 40
			        6232 => x"00000000",		-- colors: 40, 40, 40, 40
			        6233 => x"00000000",		-- colors: 40, 40, 40, 40
			        6234 => x"00000000",		-- colors: 40, 40, 40, 40
			        6235 => x"00000000",		-- colors: 40, 40, 40, 40
			        6236 => x"00000000",		-- colors: 40, 40, 40, 40
			        6237 => x"00000000",		-- colors: 40, 40, 40, 40
			        6238 => x"00000000",		-- colors: 40, 40, 40, 40
			        6239 => x"00000000",		-- colors: 40, 40, 40, 40
			        6240 => x"00000000",		-- colors: 40, 40, 40, 40
			        6241 => x"00000000",		-- colors: 40, 40, 40, 40
			        6242 => x"00000000",		-- colors: 40, 40, 40, 40
			        6243 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6244 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6245 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6246 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6247 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6248 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6249 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6250 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6251 => x"00000000",		-- colors: 40, 40, 40, 40
			        6252 => x"00000000",		-- colors: 40, 40, 40, 40
			        6253 => x"00000000",		-- colors: 40, 40, 40, 40
			        6254 => x"00000000",		-- colors: 40, 40, 40, 40
			        6255 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6256 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6257 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6258 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6259 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6260 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6261 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6262 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6263 => x"00000000",		-- colors: 40, 40, 40, 40
			        6264 => x"00000000",		-- colors: 40, 40, 40, 40
			        6265 => x"00000000",		-- colors: 40, 40, 40, 40
			        6266 => x"00000000",		-- colors: 40, 40, 40, 40
			        6267 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6268 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6269 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6270 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60

			                --  sprite 94
			        6271 => x"00000000",		-- colors: 40, 40, 40, 40
			        6272 => x"00000000",		-- colors: 40, 40, 40, 40
			        6273 => x"00000000",		-- colors: 40, 40, 40, 40
			        6274 => x"00000000",		-- colors: 40, 40, 40, 40
			        6275 => x"00000000",		-- colors: 40, 40, 40, 40
			        6276 => x"00000000",		-- colors: 40, 40, 40, 40
			        6277 => x"00000000",		-- colors: 40, 40, 40, 40
			        6278 => x"00000000",		-- colors: 40, 40, 40, 40
			        6279 => x"32323232",		-- colors: 50, 50, 50, 50
			        6280 => x"32323232",		-- colors: 50, 50, 50, 50
			        6281 => x"32323232",		-- colors: 50, 50, 50, 50
			        6282 => x"32323232",		-- colors: 50, 50, 50, 50
			        6283 => x"00000000",		-- colors: 40, 40, 40, 40
			        6284 => x"00000000",		-- colors: 40, 40, 40, 40
			        6285 => x"00000000",		-- colors: 40, 40, 40, 40
			        6286 => x"00000000",		-- colors: 40, 40, 40, 40
			        6287 => x"00000000",		-- colors: 40, 40, 40, 40
			        6288 => x"00000000",		-- colors: 40, 40, 40, 40
			        6289 => x"00000000",		-- colors: 40, 40, 40, 40
			        6290 => x"00000000",		-- colors: 40, 40, 40, 40
			        6291 => x"00000000",		-- colors: 40, 40, 40, 40
			        6292 => x"00000000",		-- colors: 40, 40, 40, 40
			        6293 => x"00000000",		-- colors: 40, 40, 40, 40
			        6294 => x"00000000",		-- colors: 40, 40, 40, 40
			        6295 => x"32323232",		-- colors: 50, 50, 50, 50
			        6296 => x"32323232",		-- colors: 50, 50, 50, 50
			        6297 => x"32323232",		-- colors: 50, 50, 50, 50
			        6298 => x"32323232",		-- colors: 50, 50, 50, 50
			        6299 => x"00000000",		-- colors: 40, 40, 40, 40
			        6300 => x"00000000",		-- colors: 40, 40, 40, 40
			        6301 => x"00000000",		-- colors: 40, 40, 40, 40
			        6302 => x"00000000",		-- colors: 40, 40, 40, 40
			        6303 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6304 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6305 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6306 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6307 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6308 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6309 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6310 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6311 => x"00000000",		-- colors: 40, 40, 40, 40
			        6312 => x"00000000",		-- colors: 40, 40, 40, 40
			        6313 => x"00000000",		-- colors: 40, 40, 40, 40
			        6314 => x"00000000",		-- colors: 40, 40, 40, 40
			        6315 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6316 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6317 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6318 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6319 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6320 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6321 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6322 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6323 => x"00000000",		-- colors: 40, 40, 40, 40
			        6324 => x"00000000",		-- colors: 40, 40, 40, 40
			        6325 => x"00000000",		-- colors: 40, 40, 40, 40
			        6326 => x"00000000",		-- colors: 40, 40, 40, 40
			        6327 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6328 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6329 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6330 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6331 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6332 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6333 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6334 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60

			                --  sprite 95
			        6335 => x"00000000",		-- colors: 40, 40, 40, 40
			        6336 => x"00000000",		-- colors: 40, 40, 40, 40
			        6337 => x"00000000",		-- colors: 40, 40, 40, 40
			        6338 => x"00000000",		-- colors: 40, 40, 40, 40
			        6339 => x"00000000",		-- colors: 40, 40, 40, 40
			        6340 => x"00000000",		-- colors: 40, 40, 40, 40
			        6341 => x"00000000",		-- colors: 40, 40, 40, 40
			        6342 => x"00000000",		-- colors: 40, 40, 40, 40
			        6343 => x"00000000",		-- colors: 40, 40, 40, 40
			        6344 => x"00000000",		-- colors: 40, 40, 40, 40
			        6345 => x"00000000",		-- colors: 40, 40, 40, 40
			        6346 => x"00000000",		-- colors: 40, 40, 40, 40
			        6347 => x"00000000",		-- colors: 40, 40, 40, 40
			        6348 => x"00000000",		-- colors: 40, 40, 40, 40
			        6349 => x"00000000",		-- colors: 40, 40, 40, 40
			        6350 => x"00000000",		-- colors: 40, 40, 40, 40
			        6351 => x"00000000",		-- colors: 40, 40, 40, 40
			        6352 => x"00000000",		-- colors: 40, 40, 40, 40
			        6353 => x"00000000",		-- colors: 40, 40, 40, 40
			        6354 => x"00000000",		-- colors: 40, 40, 40, 40
			        6355 => x"00000000",		-- colors: 40, 40, 40, 40
			        6356 => x"00000000",		-- colors: 40, 40, 40, 40
			        6357 => x"00000000",		-- colors: 40, 40, 40, 40
			        6358 => x"00000000",		-- colors: 40, 40, 40, 40
			        6359 => x"00000000",		-- colors: 40, 40, 40, 40
			        6360 => x"00000000",		-- colors: 40, 40, 40, 40
			        6361 => x"00000000",		-- colors: 40, 40, 40, 40
			        6362 => x"00000000",		-- colors: 40, 40, 40, 40
			        6363 => x"00000000",		-- colors: 40, 40, 40, 40
			        6364 => x"00000000",		-- colors: 40, 40, 40, 40
			        6365 => x"00000000",		-- colors: 40, 40, 40, 40
			        6366 => x"00000000",		-- colors: 40, 40, 40, 40
			        6367 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6368 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6369 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6370 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6371 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6372 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6373 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6374 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6375 => x"00000000",		-- colors: 40, 40, 40, 40
			        6376 => x"00000000",		-- colors: 40, 40, 40, 40
			        6377 => x"00000000",		-- colors: 40, 40, 40, 40
			        6378 => x"00000000",		-- colors: 40, 40, 40, 40
			        6379 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6380 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6381 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6382 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6383 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6384 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6385 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6386 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6387 => x"00000000",		-- colors: 40, 40, 40, 40
			        6388 => x"00000000",		-- colors: 40, 40, 40, 40
			        6389 => x"00000000",		-- colors: 40, 40, 40, 40
			        6390 => x"00000000",		-- colors: 40, 40, 40, 40
			        6391 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6392 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6393 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6394 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6395 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6396 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6397 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6398 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60

			                --  sprite 96
			        6399 => x"00000000",		-- colors: 40, 40, 40, 40
			        6400 => x"00000000",		-- colors: 40, 40, 40, 40
			        6401 => x"00000000",		-- colors: 40, 40, 40, 40
			        6402 => x"00000000",		-- colors: 40, 40, 40, 40
			        6403 => x"00000000",		-- colors: 40, 40, 40, 40
			        6404 => x"00000000",		-- colors: 40, 40, 40, 40
			        6405 => x"00000000",		-- colors: 40, 40, 40, 40
			        6406 => x"00000000",		-- colors: 40, 40, 40, 40
			        6407 => x"00000000",		-- colors: 40, 40, 40, 40
			        6408 => x"00000000",		-- colors: 40, 40, 40, 40
			        6409 => x"00000000",		-- colors: 40, 40, 40, 40
			        6410 => x"00000000",		-- colors: 40, 40, 40, 40
			        6411 => x"00000000",		-- colors: 40, 40, 40, 40
			        6412 => x"00000000",		-- colors: 40, 40, 40, 40
			        6413 => x"00000000",		-- colors: 40, 40, 40, 40
			        6414 => x"00000000",		-- colors: 40, 40, 40, 40
			        6415 => x"00000000",		-- colors: 40, 40, 40, 40
			        6416 => x"00000000",		-- colors: 40, 40, 40, 40
			        6417 => x"00000000",		-- colors: 40, 40, 40, 40
			        6418 => x"00000000",		-- colors: 40, 40, 40, 40
			        6419 => x"00000000",		-- colors: 40, 40, 40, 40
			        6420 => x"00000000",		-- colors: 40, 40, 40, 40
			        6421 => x"00000000",		-- colors: 40, 40, 40, 40
			        6422 => x"00000000",		-- colors: 40, 40, 40, 40
			        6423 => x"00000000",		-- colors: 40, 40, 40, 40
			        6424 => x"00000000",		-- colors: 40, 40, 40, 40
			        6425 => x"00000000",		-- colors: 40, 40, 40, 40
			        6426 => x"00000000",		-- colors: 40, 40, 40, 40
			        6427 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6428 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6429 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6430 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6431 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6432 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6433 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6434 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6435 => x"00000000",		-- colors: 40, 40, 40, 40
			        6436 => x"00000000",		-- colors: 40, 40, 40, 40
			        6437 => x"00000000",		-- colors: 40, 40, 40, 40
			        6438 => x"00000000",		-- colors: 40, 40, 40, 40
			        6439 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6440 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6441 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6442 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6443 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6444 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6445 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6446 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6447 => x"00000000",		-- colors: 40, 40, 40, 40
			        6448 => x"00000000",		-- colors: 40, 40, 40, 40
			        6449 => x"00000000",		-- colors: 40, 40, 40, 40
			        6450 => x"00000000",		-- colors: 40, 40, 40, 40
			        6451 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6452 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6453 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6454 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6455 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6456 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6457 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6458 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6459 => x"00000000",		-- colors: 40, 40, 40, 40
			        6460 => x"00000000",		-- colors: 40, 40, 40, 40
			        6461 => x"00000000",		-- colors: 40, 40, 40, 40
			        6462 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 97
			        6463 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6464 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6465 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6466 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6467 => x"00000000",		-- colors: 40, 40, 40, 40
			        6468 => x"00000000",		-- colors: 40, 40, 40, 40
			        6469 => x"00000000",		-- colors: 40, 40, 40, 40
			        6470 => x"00000000",		-- colors: 40, 40, 40, 40
			        6471 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6472 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6473 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6474 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6475 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6476 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6477 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6478 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6479 => x"00000000",		-- colors: 40, 40, 40, 40
			        6480 => x"00000000",		-- colors: 40, 40, 40, 40
			        6481 => x"00000000",		-- colors: 40, 40, 40, 40
			        6482 => x"00000000",		-- colors: 40, 40, 40, 40
			        6483 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6484 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6485 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6486 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6487 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6488 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6489 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6490 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6491 => x"00000000",		-- colors: 40, 40, 40, 40
			        6492 => x"00000000",		-- colors: 40, 40, 40, 40
			        6493 => x"00000000",		-- colors: 40, 40, 40, 40
			        6494 => x"00000000",		-- colors: 40, 40, 40, 40
			        6495 => x"00000000",		-- colors: 40, 40, 40, 40
			        6496 => x"00000000",		-- colors: 40, 40, 40, 40
			        6497 => x"00000000",		-- colors: 40, 40, 40, 40
			        6498 => x"00000000",		-- colors: 40, 40, 40, 40
			        6499 => x"00000000",		-- colors: 40, 40, 40, 40
			        6500 => x"00000000",		-- colors: 40, 40, 40, 40
			        6501 => x"00000000",		-- colors: 40, 40, 40, 40
			        6502 => x"00000000",		-- colors: 40, 40, 40, 40
			        6503 => x"00000000",		-- colors: 40, 40, 40, 40
			        6504 => x"00000000",		-- colors: 40, 40, 40, 40
			        6505 => x"00000000",		-- colors: 40, 40, 40, 40
			        6506 => x"00000000",		-- colors: 40, 40, 40, 40
			        6507 => x"00000000",		-- colors: 40, 40, 40, 40
			        6508 => x"00000000",		-- colors: 40, 40, 40, 40
			        6509 => x"00000000",		-- colors: 40, 40, 40, 40
			        6510 => x"00000000",		-- colors: 40, 40, 40, 40
			        6511 => x"00000000",		-- colors: 40, 40, 40, 40
			        6512 => x"00000000",		-- colors: 40, 40, 40, 40
			        6513 => x"00000000",		-- colors: 40, 40, 40, 40
			        6514 => x"00000000",		-- colors: 40, 40, 40, 40
			        6515 => x"00000000",		-- colors: 40, 40, 40, 40
			        6516 => x"00000000",		-- colors: 40, 40, 40, 40
			        6517 => x"00000000",		-- colors: 40, 40, 40, 40
			        6518 => x"00000000",		-- colors: 40, 40, 40, 40
			        6519 => x"00000000",		-- colors: 40, 40, 40, 40
			        6520 => x"00000000",		-- colors: 40, 40, 40, 40
			        6521 => x"00000000",		-- colors: 40, 40, 40, 40
			        6522 => x"00000000",		-- colors: 40, 40, 40, 40
			        6523 => x"00000000",		-- colors: 40, 40, 40, 40
			        6524 => x"00000000",		-- colors: 40, 40, 40, 40
			        6525 => x"00000000",		-- colors: 40, 40, 40, 40
			        6526 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 98
			        6527 => x"00000000",		-- colors: 40, 40, 40, 40
			        6528 => x"00000000",		-- colors: 40, 40, 40, 40
			        6529 => x"00000000",		-- colors: 40, 40, 40, 40
			        6530 => x"00000000",		-- colors: 40, 40, 40, 40
			        6531 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6532 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6533 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6534 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6535 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6536 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6537 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6538 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6539 => x"00000000",		-- colors: 40, 40, 40, 40
			        6540 => x"00000000",		-- colors: 40, 40, 40, 40
			        6541 => x"00000000",		-- colors: 40, 40, 40, 40
			        6542 => x"00000000",		-- colors: 40, 40, 40, 40
			        6543 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6544 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6545 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6546 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6547 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6548 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6549 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6550 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6551 => x"00000000",		-- colors: 40, 40, 40, 40
			        6552 => x"00000000",		-- colors: 40, 40, 40, 40
			        6553 => x"00000000",		-- colors: 40, 40, 40, 40
			        6554 => x"00000000",		-- colors: 40, 40, 40, 40
			        6555 => x"00000000",		-- colors: 40, 40, 40, 40
			        6556 => x"00000000",		-- colors: 40, 40, 40, 40
			        6557 => x"00000000",		-- colors: 40, 40, 40, 40
			        6558 => x"00000000",		-- colors: 40, 40, 40, 40
			        6559 => x"00000000",		-- colors: 40, 40, 40, 40
			        6560 => x"00000000",		-- colors: 40, 40, 40, 40
			        6561 => x"00000000",		-- colors: 40, 40, 40, 40
			        6562 => x"00000000",		-- colors: 40, 40, 40, 40
			        6563 => x"00000000",		-- colors: 40, 40, 40, 40
			        6564 => x"00000000",		-- colors: 40, 40, 40, 40
			        6565 => x"00000000",		-- colors: 40, 40, 40, 40
			        6566 => x"00000000",		-- colors: 40, 40, 40, 40
			        6567 => x"00000000",		-- colors: 40, 40, 40, 40
			        6568 => x"00000000",		-- colors: 40, 40, 40, 40
			        6569 => x"00000000",		-- colors: 40, 40, 40, 40
			        6570 => x"00000000",		-- colors: 40, 40, 40, 40
			        6571 => x"00000000",		-- colors: 40, 40, 40, 40
			        6572 => x"00000000",		-- colors: 40, 40, 40, 40
			        6573 => x"00000000",		-- colors: 40, 40, 40, 40
			        6574 => x"00000000",		-- colors: 40, 40, 40, 40
			        6575 => x"00000000",		-- colors: 40, 40, 40, 40
			        6576 => x"00000000",		-- colors: 40, 40, 40, 40
			        6577 => x"00000000",		-- colors: 40, 40, 40, 40
			        6578 => x"00000000",		-- colors: 40, 40, 40, 40
			        6579 => x"00000000",		-- colors: 40, 40, 40, 40
			        6580 => x"00000000",		-- colors: 40, 40, 40, 40
			        6581 => x"00000000",		-- colors: 40, 40, 40, 40
			        6582 => x"00000000",		-- colors: 40, 40, 40, 40
			        6583 => x"00000000",		-- colors: 40, 40, 40, 40
			        6584 => x"00000000",		-- colors: 40, 40, 40, 40
			        6585 => x"00000000",		-- colors: 40, 40, 40, 40
			        6586 => x"00000000",		-- colors: 40, 40, 40, 40
			        6587 => x"00000000",		-- colors: 40, 40, 40, 40
			        6588 => x"00000000",		-- colors: 40, 40, 40, 40
			        6589 => x"00000000",		-- colors: 40, 40, 40, 40
			        6590 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 99
			        6591 => x"00000000",		-- colors: 40, 40, 40, 40
			        6592 => x"00000000",		-- colors: 40, 40, 40, 40
			        6593 => x"00000000",		-- colors: 40, 40, 40, 40
			        6594 => x"00000000",		-- colors: 40, 40, 40, 40
			        6595 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6596 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6597 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6598 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6599 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6600 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6601 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6602 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6603 => x"00000000",		-- colors: 40, 40, 40, 40
			        6604 => x"00000000",		-- colors: 40, 40, 40, 40
			        6605 => x"00000000",		-- colors: 40, 40, 40, 40
			        6606 => x"00000000",		-- colors: 40, 40, 40, 40
			        6607 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6608 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6609 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6610 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6611 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6612 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6613 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6614 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6615 => x"00000000",		-- colors: 40, 40, 40, 40
			        6616 => x"00000000",		-- colors: 40, 40, 40, 40
			        6617 => x"00000000",		-- colors: 40, 40, 40, 40
			        6618 => x"00000000",		-- colors: 40, 40, 40, 40
			        6619 => x"00000000",		-- colors: 40, 40, 40, 40
			        6620 => x"00000000",		-- colors: 40, 40, 40, 40
			        6621 => x"00000000",		-- colors: 40, 40, 40, 40
			        6622 => x"00000000",		-- colors: 40, 40, 40, 40
			        6623 => x"00000000",		-- colors: 40, 40, 40, 40
			        6624 => x"00000000",		-- colors: 40, 40, 40, 40
			        6625 => x"00000000",		-- colors: 40, 40, 40, 40
			        6626 => x"00000000",		-- colors: 40, 40, 40, 40
			        6627 => x"00000000",		-- colors: 40, 40, 40, 40
			        6628 => x"00000000",		-- colors: 40, 40, 40, 40
			        6629 => x"00000000",		-- colors: 40, 40, 40, 40
			        6630 => x"00000000",		-- colors: 40, 40, 40, 40
			        6631 => x"00000000",		-- colors: 40, 40, 40, 40
			        6632 => x"00000000",		-- colors: 40, 40, 40, 40
			        6633 => x"00000000",		-- colors: 40, 40, 40, 40
			        6634 => x"00000000",		-- colors: 40, 40, 40, 40
			        6635 => x"00000000",		-- colors: 40, 40, 40, 40
			        6636 => x"00000000",		-- colors: 40, 40, 40, 40
			        6637 => x"00000000",		-- colors: 40, 40, 40, 40
			        6638 => x"00000000",		-- colors: 40, 40, 40, 40
			        6639 => x"00000000",		-- colors: 40, 40, 40, 40
			        6640 => x"00000000",		-- colors: 40, 40, 40, 40
			        6641 => x"00000000",		-- colors: 40, 40, 40, 40
			        6642 => x"00000000",		-- colors: 40, 40, 40, 40
			        6643 => x"00000000",		-- colors: 40, 40, 40, 40
			        6644 => x"00000000",		-- colors: 40, 40, 40, 40
			        6645 => x"00000000",		-- colors: 40, 40, 40, 40
			        6646 => x"00000000",		-- colors: 40, 40, 40, 40
			        6647 => x"00000000",		-- colors: 40, 40, 40, 40
			        6648 => x"00000000",		-- colors: 40, 40, 40, 40
			        6649 => x"00000000",		-- colors: 40, 40, 40, 40
			        6650 => x"00000000",		-- colors: 40, 40, 40, 40
			        6651 => x"00000000",		-- colors: 40, 40, 40, 40
			        6652 => x"00000000",		-- colors: 40, 40, 40, 40
			        6653 => x"00000000",		-- colors: 40, 40, 40, 40
			        6654 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 100
			        6655 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6656 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6657 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6658 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6659 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6660 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6661 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6662 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6663 => x"00000000",		-- colors: 40, 40, 40, 40
			        6664 => x"00000000",		-- colors: 40, 40, 40, 40
			        6665 => x"00000000",		-- colors: 40, 40, 40, 40
			        6666 => x"00000000",		-- colors: 40, 40, 40, 40
			        6667 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6668 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6669 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6670 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6671 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6672 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6673 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6674 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6675 => x"00000000",		-- colors: 40, 40, 40, 40
			        6676 => x"00000000",		-- colors: 40, 40, 40, 40
			        6677 => x"00000000",		-- colors: 40, 40, 40, 40
			        6678 => x"00000000",		-- colors: 40, 40, 40, 40
			        6679 => x"00000000",		-- colors: 40, 40, 40, 40
			        6680 => x"00000000",		-- colors: 40, 40, 40, 40
			        6681 => x"00000000",		-- colors: 40, 40, 40, 40
			        6682 => x"00000000",		-- colors: 40, 40, 40, 40
			        6683 => x"00000000",		-- colors: 40, 40, 40, 40
			        6684 => x"00000000",		-- colors: 40, 40, 40, 40
			        6685 => x"00000000",		-- colors: 40, 40, 40, 40
			        6686 => x"00000000",		-- colors: 40, 40, 40, 40
			        6687 => x"00000000",		-- colors: 40, 40, 40, 40
			        6688 => x"00000000",		-- colors: 40, 40, 40, 40
			        6689 => x"00000000",		-- colors: 40, 40, 40, 40
			        6690 => x"00000000",		-- colors: 40, 40, 40, 40
			        6691 => x"00000000",		-- colors: 40, 40, 40, 40
			        6692 => x"00000000",		-- colors: 40, 40, 40, 40
			        6693 => x"00000000",		-- colors: 40, 40, 40, 40
			        6694 => x"00000000",		-- colors: 40, 40, 40, 40
			        6695 => x"00000000",		-- colors: 40, 40, 40, 40
			        6696 => x"00000000",		-- colors: 40, 40, 40, 40
			        6697 => x"00000000",		-- colors: 40, 40, 40, 40
			        6698 => x"00000000",		-- colors: 40, 40, 40, 40
			        6699 => x"00000000",		-- colors: 40, 40, 40, 40
			        6700 => x"00000000",		-- colors: 40, 40, 40, 40
			        6701 => x"00000000",		-- colors: 40, 40, 40, 40
			        6702 => x"00000000",		-- colors: 40, 40, 40, 40
			        6703 => x"00000000",		-- colors: 40, 40, 40, 40
			        6704 => x"00000000",		-- colors: 40, 40, 40, 40
			        6705 => x"00000000",		-- colors: 40, 40, 40, 40
			        6706 => x"00000000",		-- colors: 40, 40, 40, 40
			        6707 => x"00000000",		-- colors: 40, 40, 40, 40
			        6708 => x"00000000",		-- colors: 40, 40, 40, 40
			        6709 => x"00000000",		-- colors: 40, 40, 40, 40
			        6710 => x"00000000",		-- colors: 40, 40, 40, 40
			        6711 => x"00000000",		-- colors: 40, 40, 40, 40
			        6712 => x"00000000",		-- colors: 40, 40, 40, 40
			        6713 => x"00000000",		-- colors: 40, 40, 40, 40
			        6714 => x"00000000",		-- colors: 40, 40, 40, 40
			        6715 => x"00000000",		-- colors: 40, 40, 40, 40
			        6716 => x"00000000",		-- colors: 40, 40, 40, 40
			        6717 => x"00000000",		-- colors: 40, 40, 40, 40
			        6718 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 101
			        6719 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6720 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6721 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6722 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6723 => x"00000000",		-- colors: 40, 40, 40, 40
			        6724 => x"00000000",		-- colors: 40, 40, 40, 40
			        6725 => x"00000000",		-- colors: 40, 40, 40, 40
			        6726 => x"00000000",		-- colors: 40, 40, 40, 40
			        6727 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6728 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6729 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6730 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6731 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6732 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6733 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6734 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6735 => x"00000000",		-- colors: 40, 40, 40, 40
			        6736 => x"00000000",		-- colors: 40, 40, 40, 40
			        6737 => x"00000000",		-- colors: 40, 40, 40, 40
			        6738 => x"00000000",		-- colors: 40, 40, 40, 40
			        6739 => x"00000000",		-- colors: 40, 40, 40, 40
			        6740 => x"00000000",		-- colors: 40, 40, 40, 40
			        6741 => x"00000000",		-- colors: 40, 40, 40, 40
			        6742 => x"00000000",		-- colors: 40, 40, 40, 40
			        6743 => x"00000000",		-- colors: 40, 40, 40, 40
			        6744 => x"00000000",		-- colors: 40, 40, 40, 40
			        6745 => x"00000000",		-- colors: 40, 40, 40, 40
			        6746 => x"00000000",		-- colors: 40, 40, 40, 40
			        6747 => x"00000000",		-- colors: 40, 40, 40, 40
			        6748 => x"00000000",		-- colors: 40, 40, 40, 40
			        6749 => x"00000000",		-- colors: 40, 40, 40, 40
			        6750 => x"00000000",		-- colors: 40, 40, 40, 40
			        6751 => x"00000000",		-- colors: 40, 40, 40, 40
			        6752 => x"00000000",		-- colors: 40, 40, 40, 40
			        6753 => x"00000000",		-- colors: 40, 40, 40, 40
			        6754 => x"00000000",		-- colors: 40, 40, 40, 40
			        6755 => x"00000000",		-- colors: 40, 40, 40, 40
			        6756 => x"00000000",		-- colors: 40, 40, 40, 40
			        6757 => x"00000000",		-- colors: 40, 40, 40, 40
			        6758 => x"00000000",		-- colors: 40, 40, 40, 40
			        6759 => x"00000000",		-- colors: 40, 40, 40, 40
			        6760 => x"00000000",		-- colors: 40, 40, 40, 40
			        6761 => x"00000000",		-- colors: 40, 40, 40, 40
			        6762 => x"00000000",		-- colors: 40, 40, 40, 40
			        6763 => x"00000000",		-- colors: 40, 40, 40, 40
			        6764 => x"00000000",		-- colors: 40, 40, 40, 40
			        6765 => x"00000000",		-- colors: 40, 40, 40, 40
			        6766 => x"00000000",		-- colors: 40, 40, 40, 40
			        6767 => x"00000000",		-- colors: 40, 40, 40, 40
			        6768 => x"00000000",		-- colors: 40, 40, 40, 40
			        6769 => x"00000000",		-- colors: 40, 40, 40, 40
			        6770 => x"00000000",		-- colors: 40, 40, 40, 40
			        6771 => x"00000000",		-- colors: 40, 40, 40, 40
			        6772 => x"00000000",		-- colors: 40, 40, 40, 40
			        6773 => x"00000000",		-- colors: 40, 40, 40, 40
			        6774 => x"00000000",		-- colors: 40, 40, 40, 40
			        6775 => x"00000000",		-- colors: 40, 40, 40, 40
			        6776 => x"00000000",		-- colors: 40, 40, 40, 40
			        6777 => x"00000000",		-- colors: 40, 40, 40, 40
			        6778 => x"00000000",		-- colors: 40, 40, 40, 40
			        6779 => x"00000000",		-- colors: 40, 40, 40, 40
			        6780 => x"00000000",		-- colors: 40, 40, 40, 40
			        6781 => x"00000000",		-- colors: 40, 40, 40, 40
			        6782 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 102
			        6783 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6784 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6785 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6786 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6787 => x"00000000",		-- colors: 40, 40, 40, 40
			        6788 => x"00000000",		-- colors: 40, 40, 40, 40
			        6789 => x"00000000",		-- colors: 40, 40, 40, 40
			        6790 => x"00000000",		-- colors: 40, 40, 40, 40
			        6791 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6792 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6793 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6794 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6795 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6796 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6797 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6798 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6799 => x"00000000",		-- colors: 40, 40, 40, 40
			        6800 => x"00000000",		-- colors: 40, 40, 40, 40
			        6801 => x"00000000",		-- colors: 40, 40, 40, 40
			        6802 => x"00000000",		-- colors: 40, 40, 40, 40
			        6803 => x"00000000",		-- colors: 40, 40, 40, 40
			        6804 => x"00000000",		-- colors: 40, 40, 40, 40
			        6805 => x"00000000",		-- colors: 40, 40, 40, 40
			        6806 => x"00000000",		-- colors: 40, 40, 40, 40
			        6807 => x"00000000",		-- colors: 40, 40, 40, 40
			        6808 => x"00000000",		-- colors: 40, 40, 40, 40
			        6809 => x"00000000",		-- colors: 40, 40, 40, 40
			        6810 => x"00000000",		-- colors: 40, 40, 40, 40
			        6811 => x"00000000",		-- colors: 40, 40, 40, 40
			        6812 => x"00000000",		-- colors: 40, 40, 40, 40
			        6813 => x"00000000",		-- colors: 40, 40, 40, 40
			        6814 => x"00000000",		-- colors: 40, 40, 40, 40
			        6815 => x"00000000",		-- colors: 40, 40, 40, 40
			        6816 => x"00000000",		-- colors: 40, 40, 40, 40
			        6817 => x"00000000",		-- colors: 40, 40, 40, 40
			        6818 => x"00000000",		-- colors: 40, 40, 40, 40
			        6819 => x"00000000",		-- colors: 40, 40, 40, 40
			        6820 => x"00000000",		-- colors: 40, 40, 40, 40
			        6821 => x"00000000",		-- colors: 40, 40, 40, 40
			        6822 => x"00000000",		-- colors: 40, 40, 40, 40
			        6823 => x"00000000",		-- colors: 40, 40, 40, 40
			        6824 => x"00000000",		-- colors: 40, 40, 40, 40
			        6825 => x"00000000",		-- colors: 40, 40, 40, 40
			        6826 => x"00000000",		-- colors: 40, 40, 40, 40
			        6827 => x"00000000",		-- colors: 40, 40, 40, 40
			        6828 => x"00000000",		-- colors: 40, 40, 40, 40
			        6829 => x"00000000",		-- colors: 40, 40, 40, 40
			        6830 => x"00000000",		-- colors: 40, 40, 40, 40
			        6831 => x"00000000",		-- colors: 40, 40, 40, 40
			        6832 => x"00000000",		-- colors: 40, 40, 40, 40
			        6833 => x"00000000",		-- colors: 40, 40, 40, 40
			        6834 => x"00000000",		-- colors: 40, 40, 40, 40
			        6835 => x"00000000",		-- colors: 40, 40, 40, 40
			        6836 => x"00000000",		-- colors: 40, 40, 40, 40
			        6837 => x"00000000",		-- colors: 40, 40, 40, 40
			        6838 => x"00000000",		-- colors: 40, 40, 40, 40
			        6839 => x"00000000",		-- colors: 40, 40, 40, 40
			        6840 => x"00000000",		-- colors: 40, 40, 40, 40
			        6841 => x"00000000",		-- colors: 40, 40, 40, 40
			        6842 => x"00000000",		-- colors: 40, 40, 40, 40
			        6843 => x"00000000",		-- colors: 40, 40, 40, 40
			        6844 => x"00000000",		-- colors: 40, 40, 40, 40
			        6845 => x"00000000",		-- colors: 40, 40, 40, 40
			        6846 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 103
			        6847 => x"00000000",		-- colors: 40, 40, 40, 40
			        6848 => x"00000000",		-- colors: 40, 40, 40, 40
			        6849 => x"00000000",		-- colors: 40, 40, 40, 40
			        6850 => x"00000000",		-- colors: 40, 40, 40, 40
			        6851 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6852 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6853 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6854 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6855 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6856 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6857 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6858 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6859 => x"00000000",		-- colors: 40, 40, 40, 40
			        6860 => x"00000000",		-- colors: 40, 40, 40, 40
			        6861 => x"00000000",		-- colors: 40, 40, 40, 40
			        6862 => x"00000000",		-- colors: 40, 40, 40, 40
			        6863 => x"00000000",		-- colors: 40, 40, 40, 40
			        6864 => x"00000000",		-- colors: 40, 40, 40, 40
			        6865 => x"00000000",		-- colors: 40, 40, 40, 40
			        6866 => x"00000000",		-- colors: 40, 40, 40, 40
			        6867 => x"00000000",		-- colors: 40, 40, 40, 40
			        6868 => x"00000000",		-- colors: 40, 40, 40, 40
			        6869 => x"00000000",		-- colors: 40, 40, 40, 40
			        6870 => x"00000000",		-- colors: 40, 40, 40, 40
			        6871 => x"00000000",		-- colors: 40, 40, 40, 40
			        6872 => x"00000000",		-- colors: 40, 40, 40, 40
			        6873 => x"00000000",		-- colors: 40, 40, 40, 40
			        6874 => x"00000000",		-- colors: 40, 40, 40, 40
			        6875 => x"00000000",		-- colors: 40, 40, 40, 40
			        6876 => x"00000000",		-- colors: 40, 40, 40, 40
			        6877 => x"00000000",		-- colors: 40, 40, 40, 40
			        6878 => x"00000000",		-- colors: 40, 40, 40, 40
			        6879 => x"00000000",		-- colors: 40, 40, 40, 40
			        6880 => x"00000000",		-- colors: 40, 40, 40, 40
			        6881 => x"00000000",		-- colors: 40, 40, 40, 40
			        6882 => x"00000000",		-- colors: 40, 40, 40, 40
			        6883 => x"00000000",		-- colors: 40, 40, 40, 40
			        6884 => x"00000000",		-- colors: 40, 40, 40, 40
			        6885 => x"00000000",		-- colors: 40, 40, 40, 40
			        6886 => x"00000000",		-- colors: 40, 40, 40, 40
			        6887 => x"00000000",		-- colors: 40, 40, 40, 40
			        6888 => x"00000000",		-- colors: 40, 40, 40, 40
			        6889 => x"00000000",		-- colors: 40, 40, 40, 40
			        6890 => x"00000000",		-- colors: 40, 40, 40, 40
			        6891 => x"00000000",		-- colors: 40, 40, 40, 40
			        6892 => x"00000000",		-- colors: 40, 40, 40, 40
			        6893 => x"00000000",		-- colors: 40, 40, 40, 40
			        6894 => x"00000000",		-- colors: 40, 40, 40, 40
			        6895 => x"00000000",		-- colors: 40, 40, 40, 40
			        6896 => x"00000000",		-- colors: 40, 40, 40, 40
			        6897 => x"00000000",		-- colors: 40, 40, 40, 40
			        6898 => x"00000000",		-- colors: 40, 40, 40, 40
			        6899 => x"00000000",		-- colors: 40, 40, 40, 40
			        6900 => x"00000000",		-- colors: 40, 40, 40, 40
			        6901 => x"00000000",		-- colors: 40, 40, 40, 40
			        6902 => x"00000000",		-- colors: 40, 40, 40, 40
			        6903 => x"00000000",		-- colors: 40, 40, 40, 40
			        6904 => x"00000000",		-- colors: 40, 40, 40, 40
			        6905 => x"00000000",		-- colors: 40, 40, 40, 40
			        6906 => x"00000000",		-- colors: 40, 40, 40, 40
			        6907 => x"00000000",		-- colors: 40, 40, 40, 40
			        6908 => x"00000000",		-- colors: 40, 40, 40, 40
			        6909 => x"00000000",		-- colors: 40, 40, 40, 40
			        6910 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 104
			        6911 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6912 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6913 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6914 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6915 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6916 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6917 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6918 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6919 => x"00000000",		-- colors: 40, 40, 40, 40
			        6920 => x"00000000",		-- colors: 40, 40, 40, 40
			        6921 => x"00000000",		-- colors: 40, 40, 40, 40
			        6922 => x"00000000",		-- colors: 40, 40, 40, 40
			        6923 => x"00000000",		-- colors: 40, 40, 40, 40
			        6924 => x"00000000",		-- colors: 40, 40, 40, 40
			        6925 => x"00000000",		-- colors: 40, 40, 40, 40
			        6926 => x"00000000",		-- colors: 40, 40, 40, 40
			        6927 => x"00000000",		-- colors: 40, 40, 40, 40
			        6928 => x"00000000",		-- colors: 40, 40, 40, 40
			        6929 => x"00000000",		-- colors: 40, 40, 40, 40
			        6930 => x"00000000",		-- colors: 40, 40, 40, 40
			        6931 => x"00000000",		-- colors: 40, 40, 40, 40
			        6932 => x"00000000",		-- colors: 40, 40, 40, 40
			        6933 => x"00000000",		-- colors: 40, 40, 40, 40
			        6934 => x"00000000",		-- colors: 40, 40, 40, 40
			        6935 => x"00000000",		-- colors: 40, 40, 40, 40
			        6936 => x"00000000",		-- colors: 40, 40, 40, 40
			        6937 => x"00000000",		-- colors: 40, 40, 40, 40
			        6938 => x"00000000",		-- colors: 40, 40, 40, 40
			        6939 => x"00000000",		-- colors: 40, 40, 40, 40
			        6940 => x"00000000",		-- colors: 40, 40, 40, 40
			        6941 => x"00000000",		-- colors: 40, 40, 40, 40
			        6942 => x"00000000",		-- colors: 40, 40, 40, 40
			        6943 => x"00000000",		-- colors: 40, 40, 40, 40
			        6944 => x"00000000",		-- colors: 40, 40, 40, 40
			        6945 => x"00000000",		-- colors: 40, 40, 40, 40
			        6946 => x"00000000",		-- colors: 40, 40, 40, 40
			        6947 => x"00000000",		-- colors: 40, 40, 40, 40
			        6948 => x"00000000",		-- colors: 40, 40, 40, 40
			        6949 => x"00000000",		-- colors: 40, 40, 40, 40
			        6950 => x"00000000",		-- colors: 40, 40, 40, 40
			        6951 => x"00000000",		-- colors: 40, 40, 40, 40
			        6952 => x"00000000",		-- colors: 40, 40, 40, 40
			        6953 => x"00000000",		-- colors: 40, 40, 40, 40
			        6954 => x"00000000",		-- colors: 40, 40, 40, 40
			        6955 => x"00000000",		-- colors: 40, 40, 40, 40
			        6956 => x"00000000",		-- colors: 40, 40, 40, 40
			        6957 => x"00000000",		-- colors: 40, 40, 40, 40
			        6958 => x"00000000",		-- colors: 40, 40, 40, 40
			        6959 => x"00000000",		-- colors: 40, 40, 40, 40
			        6960 => x"00000000",		-- colors: 40, 40, 40, 40
			        6961 => x"00000000",		-- colors: 40, 40, 40, 40
			        6962 => x"00000000",		-- colors: 40, 40, 40, 40
			        6963 => x"00000000",		-- colors: 40, 40, 40, 40
			        6964 => x"00000000",		-- colors: 40, 40, 40, 40
			        6965 => x"00000000",		-- colors: 40, 40, 40, 40
			        6966 => x"00000000",		-- colors: 40, 40, 40, 40
			        6967 => x"00000000",		-- colors: 40, 40, 40, 40
			        6968 => x"00000000",		-- colors: 40, 40, 40, 40
			        6969 => x"00000000",		-- colors: 40, 40, 40, 40
			        6970 => x"00000000",		-- colors: 40, 40, 40, 40
			        6971 => x"00000000",		-- colors: 40, 40, 40, 40
			        6972 => x"00000000",		-- colors: 40, 40, 40, 40
			        6973 => x"00000000",		-- colors: 40, 40, 40, 40
			        6974 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 105
			        6975 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6976 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6977 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6978 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6979 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6980 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6981 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6982 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        6983 => x"00000000",		-- colors: 40, 40, 40, 40
			        6984 => x"00000000",		-- colors: 40, 40, 40, 40
			        6985 => x"00000000",		-- colors: 40, 40, 40, 40
			        6986 => x"00000000",		-- colors: 40, 40, 40, 40
			        6987 => x"00000000",		-- colors: 40, 40, 40, 40
			        6988 => x"00000000",		-- colors: 40, 40, 40, 40
			        6989 => x"00000000",		-- colors: 40, 40, 40, 40
			        6990 => x"00000000",		-- colors: 40, 40, 40, 40
			        6991 => x"00000000",		-- colors: 40, 40, 40, 40
			        6992 => x"00000000",		-- colors: 40, 40, 40, 40
			        6993 => x"00000000",		-- colors: 40, 40, 40, 40
			        6994 => x"00000000",		-- colors: 40, 40, 40, 40
			        6995 => x"00000000",		-- colors: 40, 40, 40, 40
			        6996 => x"00000000",		-- colors: 40, 40, 40, 40
			        6997 => x"00000000",		-- colors: 40, 40, 40, 40
			        6998 => x"00000000",		-- colors: 40, 40, 40, 40
			        6999 => x"00000000",		-- colors: 40, 40, 40, 40
			        7000 => x"00000000",		-- colors: 40, 40, 40, 40
			        7001 => x"00000000",		-- colors: 40, 40, 40, 40
			        7002 => x"00000000",		-- colors: 40, 40, 40, 40
			        7003 => x"00000000",		-- colors: 40, 40, 40, 40
			        7004 => x"00000000",		-- colors: 40, 40, 40, 40
			        7005 => x"00000000",		-- colors: 40, 40, 40, 40
			        7006 => x"00000000",		-- colors: 40, 40, 40, 40
			        7007 => x"00000000",		-- colors: 40, 40, 40, 40
			        7008 => x"00000000",		-- colors: 40, 40, 40, 40
			        7009 => x"00000000",		-- colors: 40, 40, 40, 40
			        7010 => x"00000000",		-- colors: 40, 40, 40, 40
			        7011 => x"00000000",		-- colors: 40, 40, 40, 40
			        7012 => x"00000000",		-- colors: 40, 40, 40, 40
			        7013 => x"00000000",		-- colors: 40, 40, 40, 40
			        7014 => x"00000000",		-- colors: 40, 40, 40, 40
			        7015 => x"00000000",		-- colors: 40, 40, 40, 40
			        7016 => x"00000000",		-- colors: 40, 40, 40, 40
			        7017 => x"00000000",		-- colors: 40, 40, 40, 40
			        7018 => x"00000000",		-- colors: 40, 40, 40, 40
			        7019 => x"00000000",		-- colors: 40, 40, 40, 40
			        7020 => x"00000000",		-- colors: 40, 40, 40, 40
			        7021 => x"00000000",		-- colors: 40, 40, 40, 40
			        7022 => x"00000000",		-- colors: 40, 40, 40, 40
			        7023 => x"00000000",		-- colors: 40, 40, 40, 40
			        7024 => x"00000000",		-- colors: 40, 40, 40, 40
			        7025 => x"00000000",		-- colors: 40, 40, 40, 40
			        7026 => x"00000000",		-- colors: 40, 40, 40, 40
			        7027 => x"00000000",		-- colors: 40, 40, 40, 40
			        7028 => x"00000000",		-- colors: 40, 40, 40, 40
			        7029 => x"00000000",		-- colors: 40, 40, 40, 40
			        7030 => x"00000000",		-- colors: 40, 40, 40, 40
			        7031 => x"00000000",		-- colors: 40, 40, 40, 40
			        7032 => x"00000000",		-- colors: 40, 40, 40, 40
			        7033 => x"00000000",		-- colors: 40, 40, 40, 40
			        7034 => x"00000000",		-- colors: 40, 40, 40, 40
			        7035 => x"00000000",		-- colors: 40, 40, 40, 40
			        7036 => x"00000000",		-- colors: 40, 40, 40, 40
			        7037 => x"00000000",		-- colors: 40, 40, 40, 40
			        7038 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 106
			        7039 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7040 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7041 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7042 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7043 => x"00000000",		-- colors: 40, 40, 40, 40
			        7044 => x"00000000",		-- colors: 40, 40, 40, 40
			        7045 => x"00000000",		-- colors: 40, 40, 40, 40
			        7046 => x"00000000",		-- colors: 40, 40, 40, 40
			        7047 => x"00000000",		-- colors: 40, 40, 40, 40
			        7048 => x"00000000",		-- colors: 40, 40, 40, 40
			        7049 => x"00000000",		-- colors: 40, 40, 40, 40
			        7050 => x"00000000",		-- colors: 40, 40, 40, 40
			        7051 => x"00000000",		-- colors: 40, 40, 40, 40
			        7052 => x"00000000",		-- colors: 40, 40, 40, 40
			        7053 => x"00000000",		-- colors: 40, 40, 40, 40
			        7054 => x"00000000",		-- colors: 40, 40, 40, 40
			        7055 => x"00000000",		-- colors: 40, 40, 40, 40
			        7056 => x"00000000",		-- colors: 40, 40, 40, 40
			        7057 => x"00000000",		-- colors: 40, 40, 40, 40
			        7058 => x"00000000",		-- colors: 40, 40, 40, 40
			        7059 => x"00000000",		-- colors: 40, 40, 40, 40
			        7060 => x"00000000",		-- colors: 40, 40, 40, 40
			        7061 => x"00000000",		-- colors: 40, 40, 40, 40
			        7062 => x"00000000",		-- colors: 40, 40, 40, 40
			        7063 => x"00000000",		-- colors: 40, 40, 40, 40
			        7064 => x"00000000",		-- colors: 40, 40, 40, 40
			        7065 => x"00000000",		-- colors: 40, 40, 40, 40
			        7066 => x"00000000",		-- colors: 40, 40, 40, 40
			        7067 => x"00000000",		-- colors: 40, 40, 40, 40
			        7068 => x"00000000",		-- colors: 40, 40, 40, 40
			        7069 => x"00000000",		-- colors: 40, 40, 40, 40
			        7070 => x"00000000",		-- colors: 40, 40, 40, 40
			        7071 => x"00000000",		-- colors: 40, 40, 40, 40
			        7072 => x"00000000",		-- colors: 40, 40, 40, 40
			        7073 => x"00000000",		-- colors: 40, 40, 40, 40
			        7074 => x"00000000",		-- colors: 40, 40, 40, 40
			        7075 => x"00000000",		-- colors: 40, 40, 40, 40
			        7076 => x"00000000",		-- colors: 40, 40, 40, 40
			        7077 => x"00000000",		-- colors: 40, 40, 40, 40
			        7078 => x"00000000",		-- colors: 40, 40, 40, 40
			        7079 => x"00000000",		-- colors: 40, 40, 40, 40
			        7080 => x"00000000",		-- colors: 40, 40, 40, 40
			        7081 => x"00000000",		-- colors: 40, 40, 40, 40
			        7082 => x"00000000",		-- colors: 40, 40, 40, 40
			        7083 => x"00000000",		-- colors: 40, 40, 40, 40
			        7084 => x"00000000",		-- colors: 40, 40, 40, 40
			        7085 => x"00000000",		-- colors: 40, 40, 40, 40
			        7086 => x"00000000",		-- colors: 40, 40, 40, 40
			        7087 => x"00000000",		-- colors: 40, 40, 40, 40
			        7088 => x"00000000",		-- colors: 40, 40, 40, 40
			        7089 => x"00000000",		-- colors: 40, 40, 40, 40
			        7090 => x"00000000",		-- colors: 40, 40, 40, 40
			        7091 => x"00000000",		-- colors: 40, 40, 40, 40
			        7092 => x"00000000",		-- colors: 40, 40, 40, 40
			        7093 => x"00000000",		-- colors: 40, 40, 40, 40
			        7094 => x"00000000",		-- colors: 40, 40, 40, 40
			        7095 => x"00000000",		-- colors: 40, 40, 40, 40
			        7096 => x"00000000",		-- colors: 40, 40, 40, 40
			        7097 => x"00000000",		-- colors: 40, 40, 40, 40
			        7098 => x"00000000",		-- colors: 40, 40, 40, 40
			        7099 => x"00000000",		-- colors: 40, 40, 40, 40
			        7100 => x"00000000",		-- colors: 40, 40, 40, 40
			        7101 => x"00000000",		-- colors: 40, 40, 40, 40
			        7102 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 107
			        7103 => x"00000000",		-- colors: 40, 40, 40, 40
			        7104 => x"00000000",		-- colors: 40, 40, 40, 40
			        7105 => x"00000000",		-- colors: 40, 40, 40, 40
			        7106 => x"00000000",		-- colors: 40, 40, 40, 40
			        7107 => x"00000000",		-- colors: 40, 40, 40, 40
			        7108 => x"00000000",		-- colors: 40, 40, 40, 40
			        7109 => x"00000000",		-- colors: 40, 40, 40, 40
			        7110 => x"00000000",		-- colors: 40, 40, 40, 40
			        7111 => x"00000000",		-- colors: 40, 40, 40, 40
			        7112 => x"00000000",		-- colors: 40, 40, 40, 40
			        7113 => x"00000000",		-- colors: 40, 40, 40, 40
			        7114 => x"00000000",		-- colors: 40, 40, 40, 40
			        7115 => x"00000000",		-- colors: 40, 40, 40, 40
			        7116 => x"00000000",		-- colors: 40, 40, 40, 40
			        7117 => x"00000000",		-- colors: 40, 40, 40, 40
			        7118 => x"00000000",		-- colors: 40, 40, 40, 40
			        7119 => x"00000000",		-- colors: 40, 40, 40, 40
			        7120 => x"00000000",		-- colors: 40, 40, 40, 40
			        7121 => x"00000000",		-- colors: 40, 40, 40, 40
			        7122 => x"00000000",		-- colors: 40, 40, 40, 40
			        7123 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7124 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7125 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7126 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7127 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7128 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7129 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7130 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7131 => x"00000000",		-- colors: 40, 40, 40, 40
			        7132 => x"00000000",		-- colors: 40, 40, 40, 40
			        7133 => x"00000000",		-- colors: 40, 40, 40, 40
			        7134 => x"00000000",		-- colors: 40, 40, 40, 40
			        7135 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7136 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7137 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7138 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7139 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7140 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7141 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7142 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7143 => x"00000000",		-- colors: 40, 40, 40, 40
			        7144 => x"00000000",		-- colors: 40, 40, 40, 40
			        7145 => x"00000000",		-- colors: 40, 40, 40, 40
			        7146 => x"00000000",		-- colors: 40, 40, 40, 40
			        7147 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7148 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7149 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7150 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7151 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7152 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7153 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7154 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7155 => x"00000000",		-- colors: 40, 40, 40, 40
			        7156 => x"00000000",		-- colors: 40, 40, 40, 40
			        7157 => x"00000000",		-- colors: 40, 40, 40, 40
			        7158 => x"00000000",		-- colors: 40, 40, 40, 40
			        7159 => x"00000000",		-- colors: 40, 40, 40, 40
			        7160 => x"00000000",		-- colors: 40, 40, 40, 40
			        7161 => x"00000000",		-- colors: 40, 40, 40, 40
			        7162 => x"00000000",		-- colors: 40, 40, 40, 40
			        7163 => x"00000000",		-- colors: 40, 40, 40, 40
			        7164 => x"00000000",		-- colors: 40, 40, 40, 40
			        7165 => x"00000000",		-- colors: 40, 40, 40, 40
			        7166 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 108
			        7167 => x"00000000",		-- colors: 40, 40, 40, 40
			        7168 => x"00000000",		-- colors: 40, 40, 40, 40
			        7169 => x"00000000",		-- colors: 40, 40, 40, 40
			        7170 => x"00000000",		-- colors: 40, 40, 40, 40
			        7171 => x"00000000",		-- colors: 40, 40, 40, 40
			        7172 => x"00000000",		-- colors: 40, 40, 40, 40
			        7173 => x"00000000",		-- colors: 40, 40, 40, 40
			        7174 => x"00000000",		-- colors: 40, 40, 40, 40
			        7175 => x"00000000",		-- colors: 40, 40, 40, 40
			        7176 => x"00000000",		-- colors: 40, 40, 40, 40
			        7177 => x"00000000",		-- colors: 40, 40, 40, 40
			        7178 => x"00000000",		-- colors: 40, 40, 40, 40
			        7179 => x"00000000",		-- colors: 40, 40, 40, 40
			        7180 => x"00000000",		-- colors: 40, 40, 40, 40
			        7181 => x"00000000",		-- colors: 40, 40, 40, 40
			        7182 => x"00000000",		-- colors: 40, 40, 40, 40
			        7183 => x"00000000",		-- colors: 40, 40, 40, 40
			        7184 => x"00000000",		-- colors: 40, 40, 40, 40
			        7185 => x"00000000",		-- colors: 40, 40, 40, 40
			        7186 => x"00000000",		-- colors: 40, 40, 40, 40
			        7187 => x"00000000",		-- colors: 40, 40, 40, 40
			        7188 => x"00000000",		-- colors: 40, 40, 40, 40
			        7189 => x"00000000",		-- colors: 40, 40, 40, 40
			        7190 => x"00000000",		-- colors: 40, 40, 40, 40
			        7191 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7192 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7193 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7194 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7195 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7196 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7197 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7198 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7199 => x"00000000",		-- colors: 40, 40, 40, 40
			        7200 => x"00000000",		-- colors: 40, 40, 40, 40
			        7201 => x"00000000",		-- colors: 40, 40, 40, 40
			        7202 => x"00000000",		-- colors: 40, 40, 40, 40
			        7203 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7204 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7205 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7206 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7207 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7208 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7209 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7210 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7211 => x"00000000",		-- colors: 40, 40, 40, 40
			        7212 => x"00000000",		-- colors: 40, 40, 40, 40
			        7213 => x"00000000",		-- colors: 40, 40, 40, 40
			        7214 => x"00000000",		-- colors: 40, 40, 40, 40
			        7215 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7216 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7217 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7218 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7219 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7220 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7221 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7222 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7223 => x"00000000",		-- colors: 40, 40, 40, 40
			        7224 => x"00000000",		-- colors: 40, 40, 40, 40
			        7225 => x"00000000",		-- colors: 40, 40, 40, 40
			        7226 => x"00000000",		-- colors: 40, 40, 40, 40
			        7227 => x"00000000",		-- colors: 40, 40, 40, 40
			        7228 => x"00000000",		-- colors: 40, 40, 40, 40
			        7229 => x"00000000",		-- colors: 40, 40, 40, 40
			        7230 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 109
			        7231 => x"00000000",		-- colors: 40, 40, 40, 40
			        7232 => x"00000000",		-- colors: 40, 40, 40, 40
			        7233 => x"00000000",		-- colors: 40, 40, 40, 40
			        7234 => x"00000000",		-- colors: 40, 40, 40, 40
			        7235 => x"00000000",		-- colors: 40, 40, 40, 40
			        7236 => x"00000000",		-- colors: 40, 40, 40, 40
			        7237 => x"00000000",		-- colors: 40, 40, 40, 40
			        7238 => x"00000000",		-- colors: 40, 40, 40, 40
			        7239 => x"00000000",		-- colors: 40, 40, 40, 40
			        7240 => x"00000000",		-- colors: 40, 40, 40, 40
			        7241 => x"00000000",		-- colors: 40, 40, 40, 40
			        7242 => x"00000000",		-- colors: 40, 40, 40, 40
			        7243 => x"00000000",		-- colors: 40, 40, 40, 40
			        7244 => x"00000000",		-- colors: 40, 40, 40, 40
			        7245 => x"00000000",		-- colors: 40, 40, 40, 40
			        7246 => x"00000000",		-- colors: 40, 40, 40, 40
			        7247 => x"00000000",		-- colors: 40, 40, 40, 40
			        7248 => x"00000000",		-- colors: 40, 40, 40, 40
			        7249 => x"00000000",		-- colors: 40, 40, 40, 40
			        7250 => x"00000000",		-- colors: 40, 40, 40, 40
			        7251 => x"00000000",		-- colors: 40, 40, 40, 40
			        7252 => x"00000000",		-- colors: 40, 40, 40, 40
			        7253 => x"00000000",		-- colors: 40, 40, 40, 40
			        7254 => x"00000000",		-- colors: 40, 40, 40, 40
			        7255 => x"00000000",		-- colors: 40, 40, 40, 40
			        7256 => x"00000000",		-- colors: 40, 40, 40, 40
			        7257 => x"00000000",		-- colors: 40, 40, 40, 40
			        7258 => x"00000000",		-- colors: 40, 40, 40, 40
			        7259 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7260 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7261 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7262 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7263 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7264 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7265 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7266 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7267 => x"00000000",		-- colors: 40, 40, 40, 40
			        7268 => x"00000000",		-- colors: 40, 40, 40, 40
			        7269 => x"00000000",		-- colors: 40, 40, 40, 40
			        7270 => x"00000000",		-- colors: 40, 40, 40, 40
			        7271 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7272 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7273 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7274 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7275 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7276 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7277 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7278 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7279 => x"00000000",		-- colors: 40, 40, 40, 40
			        7280 => x"00000000",		-- colors: 40, 40, 40, 40
			        7281 => x"00000000",		-- colors: 40, 40, 40, 40
			        7282 => x"00000000",		-- colors: 40, 40, 40, 40
			        7283 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7284 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7285 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7286 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7287 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7288 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7289 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7290 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7291 => x"00000000",		-- colors: 40, 40, 40, 40
			        7292 => x"00000000",		-- colors: 40, 40, 40, 40
			        7293 => x"00000000",		-- colors: 40, 40, 40, 40
			        7294 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 110
			        7295 => x"00000000",		-- colors: 40, 40, 40, 40
			        7296 => x"00000000",		-- colors: 40, 40, 40, 40
			        7297 => x"00000000",		-- colors: 40, 40, 40, 40
			        7298 => x"00000000",		-- colors: 40, 40, 40, 40
			        7299 => x"00000000",		-- colors: 40, 40, 40, 40
			        7300 => x"00000000",		-- colors: 40, 40, 40, 40
			        7301 => x"00000000",		-- colors: 40, 40, 40, 40
			        7302 => x"00000000",		-- colors: 40, 40, 40, 40
			        7303 => x"00000000",		-- colors: 40, 40, 40, 40
			        7304 => x"00000000",		-- colors: 40, 40, 40, 40
			        7305 => x"00000000",		-- colors: 40, 40, 40, 40
			        7306 => x"00000000",		-- colors: 40, 40, 40, 40
			        7307 => x"00000000",		-- colors: 40, 40, 40, 40
			        7308 => x"00000000",		-- colors: 40, 40, 40, 40
			        7309 => x"00000000",		-- colors: 40, 40, 40, 40
			        7310 => x"00000000",		-- colors: 40, 40, 40, 40
			        7311 => x"00000000",		-- colors: 40, 40, 40, 40
			        7312 => x"00000000",		-- colors: 40, 40, 40, 40
			        7313 => x"00000000",		-- colors: 40, 40, 40, 40
			        7314 => x"00000000",		-- colors: 40, 40, 40, 40
			        7315 => x"00000000",		-- colors: 40, 40, 40, 40
			        7316 => x"00000000",		-- colors: 40, 40, 40, 40
			        7317 => x"00000000",		-- colors: 40, 40, 40, 40
			        7318 => x"00000000",		-- colors: 40, 40, 40, 40
			        7319 => x"00000000",		-- colors: 40, 40, 40, 40
			        7320 => x"00000000",		-- colors: 40, 40, 40, 40
			        7321 => x"00000000",		-- colors: 40, 40, 40, 40
			        7322 => x"00000000",		-- colors: 40, 40, 40, 40
			        7323 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7324 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7325 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7326 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7327 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7328 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7329 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7330 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7331 => x"00000000",		-- colors: 40, 40, 40, 40
			        7332 => x"00000000",		-- colors: 40, 40, 40, 40
			        7333 => x"00000000",		-- colors: 40, 40, 40, 40
			        7334 => x"00000000",		-- colors: 40, 40, 40, 40
			        7335 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7336 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7337 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7338 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7339 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7340 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7341 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7342 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7343 => x"00000000",		-- colors: 40, 40, 40, 40
			        7344 => x"00000000",		-- colors: 40, 40, 40, 40
			        7345 => x"00000000",		-- colors: 40, 40, 40, 40
			        7346 => x"00000000",		-- colors: 40, 40, 40, 40
			        7347 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7348 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7349 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7350 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7351 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7352 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7353 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7354 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7355 => x"00000000",		-- colors: 40, 40, 40, 40
			        7356 => x"00000000",		-- colors: 40, 40, 40, 40
			        7357 => x"00000000",		-- colors: 40, 40, 40, 40
			        7358 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 111
			        7359 => x"00000000",		-- colors: 40, 40, 40, 40
			        7360 => x"00000000",		-- colors: 40, 40, 40, 40
			        7361 => x"00000000",		-- colors: 40, 40, 40, 40
			        7362 => x"00000000",		-- colors: 40, 40, 40, 40
			        7363 => x"00000000",		-- colors: 40, 40, 40, 40
			        7364 => x"00000000",		-- colors: 40, 40, 40, 40
			        7365 => x"00000000",		-- colors: 40, 40, 40, 40
			        7366 => x"00000000",		-- colors: 40, 40, 40, 40
			        7367 => x"00000000",		-- colors: 40, 40, 40, 40
			        7368 => x"00000000",		-- colors: 40, 40, 40, 40
			        7369 => x"00000000",		-- colors: 40, 40, 40, 40
			        7370 => x"00000000",		-- colors: 40, 40, 40, 40
			        7371 => x"00000000",		-- colors: 40, 40, 40, 40
			        7372 => x"00000000",		-- colors: 40, 40, 40, 40
			        7373 => x"00000000",		-- colors: 40, 40, 40, 40
			        7374 => x"00000000",		-- colors: 40, 40, 40, 40
			        7375 => x"00000000",		-- colors: 40, 40, 40, 40
			        7376 => x"00000000",		-- colors: 40, 40, 40, 40
			        7377 => x"00000000",		-- colors: 40, 40, 40, 40
			        7378 => x"00000000",		-- colors: 40, 40, 40, 40
			        7379 => x"00000000",		-- colors: 40, 40, 40, 40
			        7380 => x"00000000",		-- colors: 40, 40, 40, 40
			        7381 => x"00000000",		-- colors: 40, 40, 40, 40
			        7382 => x"00000000",		-- colors: 40, 40, 40, 40
			        7383 => x"00000000",		-- colors: 40, 40, 40, 40
			        7384 => x"00000000",		-- colors: 40, 40, 40, 40
			        7385 => x"00000000",		-- colors: 40, 40, 40, 40
			        7386 => x"00000000",		-- colors: 40, 40, 40, 40
			        7387 => x"00000000",		-- colors: 40, 40, 40, 40
			        7388 => x"00000000",		-- colors: 40, 40, 40, 40
			        7389 => x"00000000",		-- colors: 40, 40, 40, 40
			        7390 => x"00000000",		-- colors: 40, 40, 40, 40
			        7391 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7392 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7393 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7394 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7395 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7396 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7397 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7398 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7399 => x"00000000",		-- colors: 40, 40, 40, 40
			        7400 => x"00000000",		-- colors: 40, 40, 40, 40
			        7401 => x"00000000",		-- colors: 40, 40, 40, 40
			        7402 => x"00000000",		-- colors: 40, 40, 40, 40
			        7403 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7404 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7405 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7406 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7407 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7408 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7409 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7410 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7411 => x"00000000",		-- colors: 40, 40, 40, 40
			        7412 => x"00000000",		-- colors: 40, 40, 40, 40
			        7413 => x"00000000",		-- colors: 40, 40, 40, 40
			        7414 => x"00000000",		-- colors: 40, 40, 40, 40
			        7415 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7416 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7417 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7418 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7419 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7420 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7421 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7422 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60

			                --  sprite 112
			        7423 => x"00000000",		-- colors: 40, 40, 40, 40
			        7424 => x"00000000",		-- colors: 40, 40, 40, 40
			        7425 => x"00000000",		-- colors: 40, 40, 40, 40
			        7426 => x"00000000",		-- colors: 40, 40, 40, 40
			        7427 => x"00000000",		-- colors: 40, 40, 40, 40
			        7428 => x"00000000",		-- colors: 40, 40, 40, 40
			        7429 => x"00000000",		-- colors: 40, 40, 40, 40
			        7430 => x"00000000",		-- colors: 40, 40, 40, 40
			        7431 => x"00000000",		-- colors: 40, 40, 40, 40
			        7432 => x"00000000",		-- colors: 40, 40, 40, 40
			        7433 => x"00000000",		-- colors: 40, 40, 40, 40
			        7434 => x"00000000",		-- colors: 40, 40, 40, 40
			        7435 => x"00000000",		-- colors: 40, 40, 40, 40
			        7436 => x"00000000",		-- colors: 40, 40, 40, 40
			        7437 => x"00000000",		-- colors: 40, 40, 40, 40
			        7438 => x"00000000",		-- colors: 40, 40, 40, 40
			        7439 => x"00000000",		-- colors: 40, 40, 40, 40
			        7440 => x"00000000",		-- colors: 40, 40, 40, 40
			        7441 => x"00000000",		-- colors: 40, 40, 40, 40
			        7442 => x"00000000",		-- colors: 40, 40, 40, 40
			        7443 => x"00000000",		-- colors: 40, 40, 40, 40
			        7444 => x"00000000",		-- colors: 40, 40, 40, 40
			        7445 => x"00000000",		-- colors: 40, 40, 40, 40
			        7446 => x"00000000",		-- colors: 40, 40, 40, 40
			        7447 => x"00000000",		-- colors: 40, 40, 40, 40
			        7448 => x"00000000",		-- colors: 40, 40, 40, 40
			        7449 => x"00000000",		-- colors: 40, 40, 40, 40
			        7450 => x"00000000",		-- colors: 40, 40, 40, 40
			        7451 => x"00000000",		-- colors: 40, 40, 40, 40
			        7452 => x"00000000",		-- colors: 40, 40, 40, 40
			        7453 => x"00000000",		-- colors: 40, 40, 40, 40
			        7454 => x"00000000",		-- colors: 40, 40, 40, 40
			        7455 => x"00000000",		-- colors: 40, 40, 40, 40
			        7456 => x"00000000",		-- colors: 40, 40, 40, 40
			        7457 => x"00000000",		-- colors: 40, 40, 40, 40
			        7458 => x"00000000",		-- colors: 40, 40, 40, 40
			        7459 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7460 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7461 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7462 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7463 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7464 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7465 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7466 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7467 => x"00000000",		-- colors: 40, 40, 40, 40
			        7468 => x"00000000",		-- colors: 40, 40, 40, 40
			        7469 => x"00000000",		-- colors: 40, 40, 40, 40
			        7470 => x"00000000",		-- colors: 40, 40, 40, 40
			        7471 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7472 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7473 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7474 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7475 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7476 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7477 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7478 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7479 => x"00000000",		-- colors: 40, 40, 40, 40
			        7480 => x"00000000",		-- colors: 40, 40, 40, 40
			        7481 => x"00000000",		-- colors: 40, 40, 40, 40
			        7482 => x"00000000",		-- colors: 40, 40, 40, 40
			        7483 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7484 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7485 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7486 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60

			                --  sprite 113
			        7487 => x"00000000",		-- colors: 40, 40, 40, 40
			        7488 => x"00000000",		-- colors: 40, 40, 40, 40
			        7489 => x"00000000",		-- colors: 40, 40, 40, 40
			        7490 => x"00000000",		-- colors: 40, 40, 40, 40
			        7491 => x"00000000",		-- colors: 40, 40, 40, 40
			        7492 => x"00000000",		-- colors: 40, 40, 40, 40
			        7493 => x"00000000",		-- colors: 40, 40, 40, 40
			        7494 => x"00000000",		-- colors: 40, 40, 40, 40
			        7495 => x"00000000",		-- colors: 40, 40, 40, 40
			        7496 => x"00000000",		-- colors: 40, 40, 40, 40
			        7497 => x"00000000",		-- colors: 40, 40, 40, 40
			        7498 => x"00000000",		-- colors: 40, 40, 40, 40
			        7499 => x"00000000",		-- colors: 40, 40, 40, 40
			        7500 => x"00000000",		-- colors: 40, 40, 40, 40
			        7501 => x"00000000",		-- colors: 40, 40, 40, 40
			        7502 => x"00000000",		-- colors: 40, 40, 40, 40
			        7503 => x"00000000",		-- colors: 40, 40, 40, 40
			        7504 => x"00000000",		-- colors: 40, 40, 40, 40
			        7505 => x"00000000",		-- colors: 40, 40, 40, 40
			        7506 => x"00000000",		-- colors: 40, 40, 40, 40
			        7507 => x"00000000",		-- colors: 40, 40, 40, 40
			        7508 => x"00000000",		-- colors: 40, 40, 40, 40
			        7509 => x"00000000",		-- colors: 40, 40, 40, 40
			        7510 => x"00000000",		-- colors: 40, 40, 40, 40
			        7511 => x"00000000",		-- colors: 40, 40, 40, 40
			        7512 => x"00000000",		-- colors: 40, 40, 40, 40
			        7513 => x"00000000",		-- colors: 40, 40, 40, 40
			        7514 => x"00000000",		-- colors: 40, 40, 40, 40
			        7515 => x"00000000",		-- colors: 40, 40, 40, 40
			        7516 => x"00000000",		-- colors: 40, 40, 40, 40
			        7517 => x"00000000",		-- colors: 40, 40, 40, 40
			        7518 => x"00000000",		-- colors: 40, 40, 40, 40
			        7519 => x"00000000",		-- colors: 40, 40, 40, 40
			        7520 => x"00000000",		-- colors: 40, 40, 40, 40
			        7521 => x"00000000",		-- colors: 40, 40, 40, 40
			        7522 => x"00000000",		-- colors: 40, 40, 40, 40
			        7523 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7524 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7525 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7526 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7527 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7528 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7529 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7530 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7531 => x"00000000",		-- colors: 40, 40, 40, 40
			        7532 => x"00000000",		-- colors: 40, 40, 40, 40
			        7533 => x"00000000",		-- colors: 40, 40, 40, 40
			        7534 => x"00000000",		-- colors: 40, 40, 40, 40
			        7535 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7536 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7537 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7538 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7539 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7540 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7541 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7542 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7543 => x"00000000",		-- colors: 40, 40, 40, 40
			        7544 => x"00000000",		-- colors: 40, 40, 40, 40
			        7545 => x"00000000",		-- colors: 40, 40, 40, 40
			        7546 => x"00000000",		-- colors: 40, 40, 40, 40
			        7547 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7548 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7549 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7550 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60

			                --  sprite 114
			        7551 => x"00000000",		-- colors: 40, 40, 40, 40
			        7552 => x"00000000",		-- colors: 40, 40, 40, 40
			        7553 => x"00000000",		-- colors: 40, 40, 40, 40
			        7554 => x"00000000",		-- colors: 40, 40, 40, 40
			        7555 => x"00000000",		-- colors: 40, 40, 40, 40
			        7556 => x"00000000",		-- colors: 40, 40, 40, 40
			        7557 => x"00000000",		-- colors: 40, 40, 40, 40
			        7558 => x"00000000",		-- colors: 40, 40, 40, 40
			        7559 => x"00000000",		-- colors: 40, 40, 40, 40
			        7560 => x"00000000",		-- colors: 40, 40, 40, 40
			        7561 => x"00000000",		-- colors: 40, 40, 40, 40
			        7562 => x"00000000",		-- colors: 40, 40, 40, 40
			        7563 => x"00000000",		-- colors: 40, 40, 40, 40
			        7564 => x"00000000",		-- colors: 40, 40, 40, 40
			        7565 => x"00000000",		-- colors: 40, 40, 40, 40
			        7566 => x"00000000",		-- colors: 40, 40, 40, 40
			        7567 => x"00000000",		-- colors: 40, 40, 40, 40
			        7568 => x"00000000",		-- colors: 40, 40, 40, 40
			        7569 => x"00000000",		-- colors: 40, 40, 40, 40
			        7570 => x"00000000",		-- colors: 40, 40, 40, 40
			        7571 => x"00000000",		-- colors: 40, 40, 40, 40
			        7572 => x"00000000",		-- colors: 40, 40, 40, 40
			        7573 => x"00000000",		-- colors: 40, 40, 40, 40
			        7574 => x"00000000",		-- colors: 40, 40, 40, 40
			        7575 => x"00000000",		-- colors: 40, 40, 40, 40
			        7576 => x"00000000",		-- colors: 40, 40, 40, 40
			        7577 => x"00000000",		-- colors: 40, 40, 40, 40
			        7578 => x"00000000",		-- colors: 40, 40, 40, 40
			        7579 => x"00000000",		-- colors: 40, 40, 40, 40
			        7580 => x"00000000",		-- colors: 40, 40, 40, 40
			        7581 => x"00000000",		-- colors: 40, 40, 40, 40
			        7582 => x"00000000",		-- colors: 40, 40, 40, 40
			        7583 => x"00000000",		-- colors: 40, 40, 40, 40
			        7584 => x"00000000",		-- colors: 40, 40, 40, 40
			        7585 => x"00000000",		-- colors: 40, 40, 40, 40
			        7586 => x"00000000",		-- colors: 40, 40, 40, 40
			        7587 => x"00000000",		-- colors: 40, 40, 40, 40
			        7588 => x"00000000",		-- colors: 40, 40, 40, 40
			        7589 => x"00000000",		-- colors: 40, 40, 40, 40
			        7590 => x"00000000",		-- colors: 40, 40, 40, 40
			        7591 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7592 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7593 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7594 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7595 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7596 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7597 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7598 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7599 => x"00000000",		-- colors: 40, 40, 40, 40
			        7600 => x"00000000",		-- colors: 40, 40, 40, 40
			        7601 => x"00000000",		-- colors: 40, 40, 40, 40
			        7602 => x"00000000",		-- colors: 40, 40, 40, 40
			        7603 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7604 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7605 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7606 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7607 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7608 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7609 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7610 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7611 => x"00000000",		-- colors: 40, 40, 40, 40
			        7612 => x"00000000",		-- colors: 40, 40, 40, 40
			        7613 => x"00000000",		-- colors: 40, 40, 40, 40
			        7614 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 115
			        7615 => x"00000000",		-- colors: 40, 40, 40, 40
			        7616 => x"00000000",		-- colors: 40, 40, 40, 40
			        7617 => x"00000000",		-- colors: 40, 40, 40, 40
			        7618 => x"00000000",		-- colors: 40, 40, 40, 40
			        7619 => x"00000000",		-- colors: 40, 40, 40, 40
			        7620 => x"00000000",		-- colors: 40, 40, 40, 40
			        7621 => x"00000000",		-- colors: 40, 40, 40, 40
			        7622 => x"00000000",		-- colors: 40, 40, 40, 40
			        7623 => x"00000000",		-- colors: 40, 40, 40, 40
			        7624 => x"00000000",		-- colors: 40, 40, 40, 40
			        7625 => x"00000000",		-- colors: 40, 40, 40, 40
			        7626 => x"00000000",		-- colors: 40, 40, 40, 40
			        7627 => x"00000000",		-- colors: 40, 40, 40, 40
			        7628 => x"00000000",		-- colors: 40, 40, 40, 40
			        7629 => x"00000000",		-- colors: 40, 40, 40, 40
			        7630 => x"00000000",		-- colors: 40, 40, 40, 40
			        7631 => x"00000000",		-- colors: 40, 40, 40, 40
			        7632 => x"00000000",		-- colors: 40, 40, 40, 40
			        7633 => x"00000000",		-- colors: 40, 40, 40, 40
			        7634 => x"00000000",		-- colors: 40, 40, 40, 40
			        7635 => x"00000000",		-- colors: 40, 40, 40, 40
			        7636 => x"00000000",		-- colors: 40, 40, 40, 40
			        7637 => x"00000000",		-- colors: 40, 40, 40, 40
			        7638 => x"00000000",		-- colors: 40, 40, 40, 40
			        7639 => x"00000000",		-- colors: 40, 40, 40, 40
			        7640 => x"00000000",		-- colors: 40, 40, 40, 40
			        7641 => x"00000000",		-- colors: 40, 40, 40, 40
			        7642 => x"00000000",		-- colors: 40, 40, 40, 40
			        7643 => x"00000000",		-- colors: 40, 40, 40, 40
			        7644 => x"00000000",		-- colors: 40, 40, 40, 40
			        7645 => x"00000000",		-- colors: 40, 40, 40, 40
			        7646 => x"00000000",		-- colors: 40, 40, 40, 40
			        7647 => x"00000000",		-- colors: 40, 40, 40, 40
			        7648 => x"00000000",		-- colors: 40, 40, 40, 40
			        7649 => x"00000000",		-- colors: 40, 40, 40, 40
			        7650 => x"00000000",		-- colors: 40, 40, 40, 40
			        7651 => x"00000000",		-- colors: 40, 40, 40, 40
			        7652 => x"00000000",		-- colors: 40, 40, 40, 40
			        7653 => x"00000000",		-- colors: 40, 40, 40, 40
			        7654 => x"00000000",		-- colors: 40, 40, 40, 40
			        7655 => x"00000000",		-- colors: 40, 40, 40, 40
			        7656 => x"00000000",		-- colors: 40, 40, 40, 40
			        7657 => x"00000000",		-- colors: 40, 40, 40, 40
			        7658 => x"00000000",		-- colors: 40, 40, 40, 40
			        7659 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7660 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7661 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7662 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7663 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7664 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7665 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7666 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7667 => x"00000000",		-- colors: 40, 40, 40, 40
			        7668 => x"00000000",		-- colors: 40, 40, 40, 40
			        7669 => x"00000000",		-- colors: 40, 40, 40, 40
			        7670 => x"00000000",		-- colors: 40, 40, 40, 40
			        7671 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7672 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7673 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7674 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7675 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7676 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7677 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7678 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60

			                --  sprite 116
			        7679 => x"00000000",		-- colors: 40, 40, 40, 40
			        7680 => x"00000000",		-- colors: 40, 40, 40, 40
			        7681 => x"00000000",		-- colors: 40, 40, 40, 40
			        7682 => x"00000000",		-- colors: 40, 40, 40, 40
			        7683 => x"00000000",		-- colors: 40, 40, 40, 40
			        7684 => x"00000000",		-- colors: 40, 40, 40, 40
			        7685 => x"00000000",		-- colors: 40, 40, 40, 40
			        7686 => x"00000000",		-- colors: 40, 40, 40, 40
			        7687 => x"00000000",		-- colors: 40, 40, 40, 40
			        7688 => x"00000000",		-- colors: 40, 40, 40, 40
			        7689 => x"00000000",		-- colors: 40, 40, 40, 40
			        7690 => x"00000000",		-- colors: 40, 40, 40, 40
			        7691 => x"00000000",		-- colors: 40, 40, 40, 40
			        7692 => x"00000000",		-- colors: 40, 40, 40, 40
			        7693 => x"00000000",		-- colors: 40, 40, 40, 40
			        7694 => x"00000000",		-- colors: 40, 40, 40, 40
			        7695 => x"00000000",		-- colors: 40, 40, 40, 40
			        7696 => x"00000000",		-- colors: 40, 40, 40, 40
			        7697 => x"00000000",		-- colors: 40, 40, 40, 40
			        7698 => x"00000000",		-- colors: 40, 40, 40, 40
			        7699 => x"00000000",		-- colors: 40, 40, 40, 40
			        7700 => x"00000000",		-- colors: 40, 40, 40, 40
			        7701 => x"00000000",		-- colors: 40, 40, 40, 40
			        7702 => x"00000000",		-- colors: 40, 40, 40, 40
			        7703 => x"00000000",		-- colors: 40, 40, 40, 40
			        7704 => x"00000000",		-- colors: 40, 40, 40, 40
			        7705 => x"00000000",		-- colors: 40, 40, 40, 40
			        7706 => x"00000000",		-- colors: 40, 40, 40, 40
			        7707 => x"00000000",		-- colors: 40, 40, 40, 40
			        7708 => x"00000000",		-- colors: 40, 40, 40, 40
			        7709 => x"00000000",		-- colors: 40, 40, 40, 40
			        7710 => x"00000000",		-- colors: 40, 40, 40, 40
			        7711 => x"00000000",		-- colors: 40, 40, 40, 40
			        7712 => x"00000000",		-- colors: 40, 40, 40, 40
			        7713 => x"00000000",		-- colors: 40, 40, 40, 40
			        7714 => x"00000000",		-- colors: 40, 40, 40, 40
			        7715 => x"00000000",		-- colors: 40, 40, 40, 40
			        7716 => x"00000000",		-- colors: 40, 40, 40, 40
			        7717 => x"00000000",		-- colors: 40, 40, 40, 40
			        7718 => x"00000000",		-- colors: 40, 40, 40, 40
			        7719 => x"00000000",		-- colors: 40, 40, 40, 40
			        7720 => x"00000000",		-- colors: 40, 40, 40, 40
			        7721 => x"00000000",		-- colors: 40, 40, 40, 40
			        7722 => x"00000000",		-- colors: 40, 40, 40, 40
			        7723 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7724 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7725 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7726 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7727 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7728 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7729 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7730 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7731 => x"00000000",		-- colors: 40, 40, 40, 40
			        7732 => x"00000000",		-- colors: 40, 40, 40, 40
			        7733 => x"00000000",		-- colors: 40, 40, 40, 40
			        7734 => x"00000000",		-- colors: 40, 40, 40, 40
			        7735 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7736 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7737 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7738 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7739 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7740 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7741 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7742 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60

			                --  sprite 117
			        7743 => x"00000000",		-- colors: 40, 40, 40, 40
			        7744 => x"00000000",		-- colors: 40, 40, 40, 40
			        7745 => x"00000000",		-- colors: 40, 40, 40, 40
			        7746 => x"00000000",		-- colors: 40, 40, 40, 40
			        7747 => x"00000000",		-- colors: 40, 40, 40, 40
			        7748 => x"00000000",		-- colors: 40, 40, 40, 40
			        7749 => x"00000000",		-- colors: 40, 40, 40, 40
			        7750 => x"00000000",		-- colors: 40, 40, 40, 40
			        7751 => x"00000000",		-- colors: 40, 40, 40, 40
			        7752 => x"00000000",		-- colors: 40, 40, 40, 40
			        7753 => x"00000000",		-- colors: 40, 40, 40, 40
			        7754 => x"00000000",		-- colors: 40, 40, 40, 40
			        7755 => x"00000000",		-- colors: 40, 40, 40, 40
			        7756 => x"00000000",		-- colors: 40, 40, 40, 40
			        7757 => x"00000000",		-- colors: 40, 40, 40, 40
			        7758 => x"00000000",		-- colors: 40, 40, 40, 40
			        7759 => x"00000000",		-- colors: 40, 40, 40, 40
			        7760 => x"00000000",		-- colors: 40, 40, 40, 40
			        7761 => x"00000000",		-- colors: 40, 40, 40, 40
			        7762 => x"00000000",		-- colors: 40, 40, 40, 40
			        7763 => x"00000000",		-- colors: 40, 40, 40, 40
			        7764 => x"00000000",		-- colors: 40, 40, 40, 40
			        7765 => x"00000000",		-- colors: 40, 40, 40, 40
			        7766 => x"00000000",		-- colors: 40, 40, 40, 40
			        7767 => x"00000000",		-- colors: 40, 40, 40, 40
			        7768 => x"00000000",		-- colors: 40, 40, 40, 40
			        7769 => x"00000000",		-- colors: 40, 40, 40, 40
			        7770 => x"00000000",		-- colors: 40, 40, 40, 40
			        7771 => x"00000000",		-- colors: 40, 40, 40, 40
			        7772 => x"00000000",		-- colors: 40, 40, 40, 40
			        7773 => x"00000000",		-- colors: 40, 40, 40, 40
			        7774 => x"00000000",		-- colors: 40, 40, 40, 40
			        7775 => x"00000000",		-- colors: 40, 40, 40, 40
			        7776 => x"00000000",		-- colors: 40, 40, 40, 40
			        7777 => x"00000000",		-- colors: 40, 40, 40, 40
			        7778 => x"00000000",		-- colors: 40, 40, 40, 40
			        7779 => x"00000000",		-- colors: 40, 40, 40, 40
			        7780 => x"00000000",		-- colors: 40, 40, 40, 40
			        7781 => x"00000000",		-- colors: 40, 40, 40, 40
			        7782 => x"00000000",		-- colors: 40, 40, 40, 40
			        7783 => x"00000000",		-- colors: 40, 40, 40, 40
			        7784 => x"00000000",		-- colors: 40, 40, 40, 40
			        7785 => x"00000000",		-- colors: 40, 40, 40, 40
			        7786 => x"00000000",		-- colors: 40, 40, 40, 40
			        7787 => x"00000000",		-- colors: 40, 40, 40, 40
			        7788 => x"00000000",		-- colors: 40, 40, 40, 40
			        7789 => x"00000000",		-- colors: 40, 40, 40, 40
			        7790 => x"00000000",		-- colors: 40, 40, 40, 40
			        7791 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7792 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7793 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7794 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7795 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7796 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7797 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7798 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7799 => x"00000000",		-- colors: 40, 40, 40, 40
			        7800 => x"00000000",		-- colors: 40, 40, 40, 40
			        7801 => x"00000000",		-- colors: 40, 40, 40, 40
			        7802 => x"00000000",		-- colors: 40, 40, 40, 40
			        7803 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7804 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7805 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7806 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60

			                --  sprite 118
			        7807 => x"00000000",		-- colors: 40, 40, 40, 40
			        7808 => x"00000000",		-- colors: 40, 40, 40, 40
			        7809 => x"00000000",		-- colors: 40, 40, 40, 40
			        7810 => x"00000000",		-- colors: 40, 40, 40, 40
			        7811 => x"00000000",		-- colors: 40, 40, 40, 40
			        7812 => x"00000000",		-- colors: 40, 40, 40, 40
			        7813 => x"00000000",		-- colors: 40, 40, 40, 40
			        7814 => x"00000000",		-- colors: 40, 40, 40, 40
			        7815 => x"00000000",		-- colors: 40, 40, 40, 40
			        7816 => x"00000000",		-- colors: 40, 40, 40, 40
			        7817 => x"00000000",		-- colors: 40, 40, 40, 40
			        7818 => x"00000000",		-- colors: 40, 40, 40, 40
			        7819 => x"00000000",		-- colors: 40, 40, 40, 40
			        7820 => x"00000000",		-- colors: 40, 40, 40, 40
			        7821 => x"00000000",		-- colors: 40, 40, 40, 40
			        7822 => x"00000000",		-- colors: 40, 40, 40, 40
			        7823 => x"00000000",		-- colors: 40, 40, 40, 40
			        7824 => x"00000000",		-- colors: 40, 40, 40, 40
			        7825 => x"00000000",		-- colors: 40, 40, 40, 40
			        7826 => x"00000000",		-- colors: 40, 40, 40, 40
			        7827 => x"00000000",		-- colors: 40, 40, 40, 40
			        7828 => x"00000000",		-- colors: 40, 40, 40, 40
			        7829 => x"00000000",		-- colors: 40, 40, 40, 40
			        7830 => x"00000000",		-- colors: 40, 40, 40, 40
			        7831 => x"00000000",		-- colors: 40, 40, 40, 40
			        7832 => x"00000000",		-- colors: 40, 40, 40, 40
			        7833 => x"00000000",		-- colors: 40, 40, 40, 40
			        7834 => x"00000000",		-- colors: 40, 40, 40, 40
			        7835 => x"00000000",		-- colors: 40, 40, 40, 40
			        7836 => x"00000000",		-- colors: 40, 40, 40, 40
			        7837 => x"00000000",		-- colors: 40, 40, 40, 40
			        7838 => x"00000000",		-- colors: 40, 40, 40, 40
			        7839 => x"00000000",		-- colors: 40, 40, 40, 40
			        7840 => x"00000000",		-- colors: 40, 40, 40, 40
			        7841 => x"00000000",		-- colors: 40, 40, 40, 40
			        7842 => x"00000000",		-- colors: 40, 40, 40, 40
			        7843 => x"00000000",		-- colors: 40, 40, 40, 40
			        7844 => x"00000000",		-- colors: 40, 40, 40, 40
			        7845 => x"00000000",		-- colors: 40, 40, 40, 40
			        7846 => x"00000000",		-- colors: 40, 40, 40, 40
			        7847 => x"00000000",		-- colors: 40, 40, 40, 40
			        7848 => x"00000000",		-- colors: 40, 40, 40, 40
			        7849 => x"00000000",		-- colors: 40, 40, 40, 40
			        7850 => x"00000000",		-- colors: 40, 40, 40, 40
			        7851 => x"00000000",		-- colors: 40, 40, 40, 40
			        7852 => x"00000000",		-- colors: 40, 40, 40, 40
			        7853 => x"00000000",		-- colors: 40, 40, 40, 40
			        7854 => x"00000000",		-- colors: 40, 40, 40, 40
			        7855 => x"00000000",		-- colors: 40, 40, 40, 40
			        7856 => x"00000000",		-- colors: 40, 40, 40, 40
			        7857 => x"00000000",		-- colors: 40, 40, 40, 40
			        7858 => x"00000000",		-- colors: 40, 40, 40, 40
			        7859 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7860 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7861 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7862 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7863 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7864 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7865 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7866 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7867 => x"00000000",		-- colors: 40, 40, 40, 40
			        7868 => x"00000000",		-- colors: 40, 40, 40, 40
			        7869 => x"00000000",		-- colors: 40, 40, 40, 40
			        7870 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 119
			        7871 => x"00000000",		-- colors: 40, 40, 40, 40
			        7872 => x"00000000",		-- colors: 40, 40, 40, 40
			        7873 => x"00000000",		-- colors: 40, 40, 40, 40
			        7874 => x"00000000",		-- colors: 40, 40, 40, 40
			        7875 => x"00000000",		-- colors: 40, 40, 40, 40
			        7876 => x"00000000",		-- colors: 40, 40, 40, 40
			        7877 => x"00000000",		-- colors: 40, 40, 40, 40
			        7878 => x"00000000",		-- colors: 40, 40, 40, 40
			        7879 => x"00000000",		-- colors: 40, 40, 40, 40
			        7880 => x"00000000",		-- colors: 40, 40, 40, 40
			        7881 => x"00000000",		-- colors: 40, 40, 40, 40
			        7882 => x"00000000",		-- colors: 40, 40, 40, 40
			        7883 => x"00000000",		-- colors: 40, 40, 40, 40
			        7884 => x"00000000",		-- colors: 40, 40, 40, 40
			        7885 => x"00000000",		-- colors: 40, 40, 40, 40
			        7886 => x"00000000",		-- colors: 40, 40, 40, 40
			        7887 => x"00000000",		-- colors: 40, 40, 40, 40
			        7888 => x"00000000",		-- colors: 40, 40, 40, 40
			        7889 => x"00000000",		-- colors: 40, 40, 40, 40
			        7890 => x"00000000",		-- colors: 40, 40, 40, 40
			        7891 => x"00000000",		-- colors: 40, 40, 40, 40
			        7892 => x"00000000",		-- colors: 40, 40, 40, 40
			        7893 => x"00000000",		-- colors: 40, 40, 40, 40
			        7894 => x"00000000",		-- colors: 40, 40, 40, 40
			        7895 => x"00000000",		-- colors: 40, 40, 40, 40
			        7896 => x"00000000",		-- colors: 40, 40, 40, 40
			        7897 => x"00000000",		-- colors: 40, 40, 40, 40
			        7898 => x"00000000",		-- colors: 40, 40, 40, 40
			        7899 => x"00000000",		-- colors: 40, 40, 40, 40
			        7900 => x"00000000",		-- colors: 40, 40, 40, 40
			        7901 => x"00000000",		-- colors: 40, 40, 40, 40
			        7902 => x"00000000",		-- colors: 40, 40, 40, 40
			        7903 => x"00000000",		-- colors: 40, 40, 40, 40
			        7904 => x"00000000",		-- colors: 40, 40, 40, 40
			        7905 => x"00000000",		-- colors: 40, 40, 40, 40
			        7906 => x"00000000",		-- colors: 40, 40, 40, 40
			        7907 => x"00000000",		-- colors: 40, 40, 40, 40
			        7908 => x"00000000",		-- colors: 40, 40, 40, 40
			        7909 => x"00000000",		-- colors: 40, 40, 40, 40
			        7910 => x"00000000",		-- colors: 40, 40, 40, 40
			        7911 => x"00000000",		-- colors: 40, 40, 40, 40
			        7912 => x"00000000",		-- colors: 40, 40, 40, 40
			        7913 => x"00000000",		-- colors: 40, 40, 40, 40
			        7914 => x"00000000",		-- colors: 40, 40, 40, 40
			        7915 => x"00000000",		-- colors: 40, 40, 40, 40
			        7916 => x"00000000",		-- colors: 40, 40, 40, 40
			        7917 => x"00000000",		-- colors: 40, 40, 40, 40
			        7918 => x"00000000",		-- colors: 40, 40, 40, 40
			        7919 => x"00000000",		-- colors: 40, 40, 40, 40
			        7920 => x"00000000",		-- colors: 40, 40, 40, 40
			        7921 => x"00000000",		-- colors: 40, 40, 40, 40
			        7922 => x"00000000",		-- colors: 40, 40, 40, 40
			        7923 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7924 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7925 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7926 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7927 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7928 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7929 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7930 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        7931 => x"00000000",		-- colors: 40, 40, 40, 40
			        7932 => x"00000000",		-- colors: 40, 40, 40, 40
			        7933 => x"00000000",		-- colors: 40, 40, 40, 40
			        7934 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 120
			        7935 => x"00000000",		-- colors: 40, 40, 40, 40
			        7936 => x"00000000",		-- colors: 40, 40, 40, 40
			        7937 => x"00000000",		-- colors: 40, 40, 40, 40
			        7938 => x"00000000",		-- colors: 40, 40, 40, 40
			        7939 => x"00000000",		-- colors: 40, 40, 40, 40
			        7940 => x"00000000",		-- colors: 40, 40, 40, 40
			        7941 => x"00000000",		-- colors: 40, 40, 40, 40
			        7942 => x"00000000",		-- colors: 40, 40, 40, 40
			        7943 => x"00000000",		-- colors: 40, 40, 40, 40
			        7944 => x"00000000",		-- colors: 40, 40, 40, 40
			        7945 => x"00000000",		-- colors: 40, 40, 40, 40
			        7946 => x"00000000",		-- colors: 40, 40, 40, 40
			        7947 => x"00000000",		-- colors: 40, 40, 40, 40
			        7948 => x"00000000",		-- colors: 40, 40, 40, 40
			        7949 => x"00000000",		-- colors: 40, 40, 40, 40
			        7950 => x"00000000",		-- colors: 40, 40, 40, 40
			        7951 => x"00000000",		-- colors: 40, 40, 40, 40
			        7952 => x"00000000",		-- colors: 40, 40, 40, 40
			        7953 => x"00000000",		-- colors: 40, 40, 40, 40
			        7954 => x"00000000",		-- colors: 40, 40, 40, 40
			        7955 => x"00000000",		-- colors: 40, 40, 40, 40
			        7956 => x"00000000",		-- colors: 40, 40, 40, 40
			        7957 => x"00000000",		-- colors: 40, 40, 40, 40
			        7958 => x"00000000",		-- colors: 40, 40, 40, 40
			        7959 => x"00000000",		-- colors: 40, 40, 40, 40
			        7960 => x"00000000",		-- colors: 40, 40, 40, 40
			        7961 => x"00000000",		-- colors: 40, 40, 40, 40
			        7962 => x"00000000",		-- colors: 40, 40, 40, 40
			        7963 => x"00000000",		-- colors: 40, 40, 40, 40
			        7964 => x"00000000",		-- colors: 40, 40, 40, 40
			        7965 => x"00000000",		-- colors: 40, 40, 40, 40
			        7966 => x"00000000",		-- colors: 40, 40, 40, 40
			        7967 => x"00000000",		-- colors: 40, 40, 40, 40
			        7968 => x"00000000",		-- colors: 40, 40, 40, 40
			        7969 => x"00000000",		-- colors: 40, 40, 40, 40
			        7970 => x"00000000",		-- colors: 40, 40, 40, 40
			        7971 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
			        7972 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
			        7973 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
			        7974 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
			        7975 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
			        7976 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
			        7977 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
			        7978 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
			        7979 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
			        7980 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
			        7981 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
			        7982 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
			        7983 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
			        7984 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
			        7985 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
			        7986 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
			        7987 => x"32323232",		-- colors: 50, 50, 50, 50
			        7988 => x"32323232",		-- colors: 50, 50, 50, 50
			        7989 => x"32323232",		-- colors: 50, 50, 50, 50
			        7990 => x"32323232",		-- colors: 50, 50, 50, 50
			        7991 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
			        7992 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
			        7993 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
			        7994 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
			        7995 => x"32323232",		-- colors: 50, 50, 50, 50
			        7996 => x"32323232",		-- colors: 50, 50, 50, 50
			        7997 => x"32323232",		-- colors: 50, 50, 50, 50
			        7998 => x"32323232",		-- colors: 50, 50, 50, 50

			                --  sprite 121
			        7999 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8000 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8001 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8002 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8003 => x"00000000",		-- colors: 40, 40, 40, 40
			        8004 => x"00000000",		-- colors: 40, 40, 40, 40
			        8005 => x"00000000",		-- colors: 40, 40, 40, 40
			        8006 => x"00000000",		-- colors: 40, 40, 40, 40
			        8007 => x"00000000",		-- colors: 40, 40, 40, 40
			        8008 => x"00000000",		-- colors: 40, 40, 40, 40
			        8009 => x"00000000",		-- colors: 40, 40, 40, 40
			        8010 => x"00000000",		-- colors: 40, 40, 40, 40
			        8011 => x"00000000",		-- colors: 40, 40, 40, 40
			        8012 => x"00000000",		-- colors: 40, 40, 40, 40
			        8013 => x"00000000",		-- colors: 40, 40, 40, 40
			        8014 => x"00000000",		-- colors: 40, 40, 40, 40
			        8015 => x"00000000",		-- colors: 40, 40, 40, 40
			        8016 => x"00000000",		-- colors: 40, 40, 40, 40
			        8017 => x"00000000",		-- colors: 40, 40, 40, 40
			        8018 => x"00000000",		-- colors: 40, 40, 40, 40
			        8019 => x"00000000",		-- colors: 40, 40, 40, 40
			        8020 => x"00000000",		-- colors: 40, 40, 40, 40
			        8021 => x"00000000",		-- colors: 40, 40, 40, 40
			        8022 => x"00000000",		-- colors: 40, 40, 40, 40
			        8023 => x"00000000",		-- colors: 40, 40, 40, 40
			        8024 => x"00000000",		-- colors: 40, 40, 40, 40
			        8025 => x"00000000",		-- colors: 40, 40, 40, 40
			        8026 => x"00000000",		-- colors: 40, 40, 40, 40
			        8027 => x"00000000",		-- colors: 40, 40, 40, 40
			        8028 => x"00000000",		-- colors: 40, 40, 40, 40
			        8029 => x"00000000",		-- colors: 40, 40, 40, 40
			        8030 => x"00000000",		-- colors: 40, 40, 40, 40
			        8031 => x"00000000",		-- colors: 40, 40, 40, 40
			        8032 => x"00000000",		-- colors: 40, 40, 40, 40
			        8033 => x"00000000",		-- colors: 40, 40, 40, 40
			        8034 => x"00000000",		-- colors: 40, 40, 40, 40
			        8035 => x"00000000",		-- colors: 40, 40, 40, 40
			        8036 => x"00000000",		-- colors: 40, 40, 40, 40
			        8037 => x"00000000",		-- colors: 40, 40, 40, 40
			        8038 => x"00000000",		-- colors: 40, 40, 40, 40
			        8039 => x"00000000",		-- colors: 40, 40, 40, 40
			        8040 => x"00000000",		-- colors: 40, 40, 40, 40
			        8041 => x"00000000",		-- colors: 40, 40, 40, 40
			        8042 => x"00000000",		-- colors: 40, 40, 40, 40
			        8043 => x"00000000",		-- colors: 40, 40, 40, 40
			        8044 => x"00000000",		-- colors: 40, 40, 40, 40
			        8045 => x"00000000",		-- colors: 40, 40, 40, 40
			        8046 => x"00000000",		-- colors: 40, 40, 40, 40
			        8047 => x"00000000",		-- colors: 40, 40, 40, 40
			        8048 => x"00000000",		-- colors: 40, 40, 40, 40
			        8049 => x"00000000",		-- colors: 40, 40, 40, 40
			        8050 => x"00000000",		-- colors: 40, 40, 40, 40
			        8051 => x"00000000",		-- colors: 40, 40, 40, 40
			        8052 => x"00000000",		-- colors: 40, 40, 40, 40
			        8053 => x"00000000",		-- colors: 40, 40, 40, 40
			        8054 => x"00000000",		-- colors: 40, 40, 40, 40
			        8055 => x"00000000",		-- colors: 40, 40, 40, 40
			        8056 => x"00000000",		-- colors: 40, 40, 40, 40
			        8057 => x"00000000",		-- colors: 40, 40, 40, 40
			        8058 => x"00000000",		-- colors: 40, 40, 40, 40
			        8059 => x"00000000",		-- colors: 40, 40, 40, 40
			        8060 => x"00000000",		-- colors: 40, 40, 40, 40
			        8061 => x"00000000",		-- colors: 40, 40, 40, 40
			        8062 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 122
			        8063 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8064 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8065 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8066 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8067 => x"00000000",		-- colors: 40, 40, 40, 40
			        8068 => x"00000000",		-- colors: 40, 40, 40, 40
			        8069 => x"00000000",		-- colors: 40, 40, 40, 40
			        8070 => x"00000000",		-- colors: 40, 40, 40, 40
			        8071 => x"00000000",		-- colors: 40, 40, 40, 40
			        8072 => x"00000000",		-- colors: 40, 40, 40, 40
			        8073 => x"00000000",		-- colors: 40, 40, 40, 40
			        8074 => x"00000000",		-- colors: 40, 40, 40, 40
			        8075 => x"00000000",		-- colors: 40, 40, 40, 40
			        8076 => x"00000000",		-- colors: 40, 40, 40, 40
			        8077 => x"00000000",		-- colors: 40, 40, 40, 40
			        8078 => x"00000000",		-- colors: 40, 40, 40, 40
			        8079 => x"00000000",		-- colors: 40, 40, 40, 40
			        8080 => x"00000000",		-- colors: 40, 40, 40, 40
			        8081 => x"00000000",		-- colors: 40, 40, 40, 40
			        8082 => x"00000000",		-- colors: 40, 40, 40, 40
			        8083 => x"00000000",		-- colors: 40, 40, 40, 40
			        8084 => x"00000000",		-- colors: 40, 40, 40, 40
			        8085 => x"00000000",		-- colors: 40, 40, 40, 40
			        8086 => x"00000000",		-- colors: 40, 40, 40, 40
			        8087 => x"00000000",		-- colors: 40, 40, 40, 40
			        8088 => x"00000000",		-- colors: 40, 40, 40, 40
			        8089 => x"00000000",		-- colors: 40, 40, 40, 40
			        8090 => x"00000000",		-- colors: 40, 40, 40, 40
			        8091 => x"00000000",		-- colors: 40, 40, 40, 40
			        8092 => x"00000000",		-- colors: 40, 40, 40, 40
			        8093 => x"00000000",		-- colors: 40, 40, 40, 40
			        8094 => x"00000000",		-- colors: 40, 40, 40, 40
			        8095 => x"00000000",		-- colors: 40, 40, 40, 40
			        8096 => x"00000000",		-- colors: 40, 40, 40, 40
			        8097 => x"00000000",		-- colors: 40, 40, 40, 40
			        8098 => x"00000000",		-- colors: 40, 40, 40, 40
			        8099 => x"00000000",		-- colors: 40, 40, 40, 40
			        8100 => x"00000000",		-- colors: 40, 40, 40, 40
			        8101 => x"00000000",		-- colors: 40, 40, 40, 40
			        8102 => x"00000000",		-- colors: 40, 40, 40, 40
			        8103 => x"00000000",		-- colors: 40, 40, 40, 40
			        8104 => x"00000000",		-- colors: 40, 40, 40, 40
			        8105 => x"00000000",		-- colors: 40, 40, 40, 40
			        8106 => x"00000000",		-- colors: 40, 40, 40, 40
			        8107 => x"00000000",		-- colors: 40, 40, 40, 40
			        8108 => x"00000000",		-- colors: 40, 40, 40, 40
			        8109 => x"00000000",		-- colors: 40, 40, 40, 40
			        8110 => x"00000000",		-- colors: 40, 40, 40, 40
			        8111 => x"00000000",		-- colors: 40, 40, 40, 40
			        8112 => x"00000000",		-- colors: 40, 40, 40, 40
			        8113 => x"00000000",		-- colors: 40, 40, 40, 40
			        8114 => x"00000000",		-- colors: 40, 40, 40, 40
			        8115 => x"00000000",		-- colors: 40, 40, 40, 40
			        8116 => x"00000000",		-- colors: 40, 40, 40, 40
			        8117 => x"00000000",		-- colors: 40, 40, 40, 40
			        8118 => x"00000000",		-- colors: 40, 40, 40, 40
			        8119 => x"00000000",		-- colors: 40, 40, 40, 40
			        8120 => x"00000000",		-- colors: 40, 40, 40, 40
			        8121 => x"00000000",		-- colors: 40, 40, 40, 40
			        8122 => x"00000000",		-- colors: 40, 40, 40, 40
			        8123 => x"00000000",		-- colors: 40, 40, 40, 40
			        8124 => x"00000000",		-- colors: 40, 40, 40, 40
			        8125 => x"00000000",		-- colors: 40, 40, 40, 40
			        8126 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 123
			        8127 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8128 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8129 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8130 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8131 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8132 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8133 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8134 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8135 => x"00000000",		-- colors: 40, 40, 40, 40
			        8136 => x"00000000",		-- colors: 40, 40, 40, 40
			        8137 => x"00000000",		-- colors: 40, 40, 40, 40
			        8138 => x"00000000",		-- colors: 40, 40, 40, 40
			        8139 => x"00000000",		-- colors: 40, 40, 40, 40
			        8140 => x"00000000",		-- colors: 40, 40, 40, 40
			        8141 => x"00000000",		-- colors: 40, 40, 40, 40
			        8142 => x"00000000",		-- colors: 40, 40, 40, 40
			        8143 => x"00000000",		-- colors: 40, 40, 40, 40
			        8144 => x"00000000",		-- colors: 40, 40, 40, 40
			        8145 => x"00000000",		-- colors: 40, 40, 40, 40
			        8146 => x"00000000",		-- colors: 40, 40, 40, 40
			        8147 => x"00000000",		-- colors: 40, 40, 40, 40
			        8148 => x"00000000",		-- colors: 40, 40, 40, 40
			        8149 => x"00000000",		-- colors: 40, 40, 40, 40
			        8150 => x"00000000",		-- colors: 40, 40, 40, 40
			        8151 => x"00000000",		-- colors: 40, 40, 40, 40
			        8152 => x"00000000",		-- colors: 40, 40, 40, 40
			        8153 => x"00000000",		-- colors: 40, 40, 40, 40
			        8154 => x"00000000",		-- colors: 40, 40, 40, 40
			        8155 => x"00000000",		-- colors: 40, 40, 40, 40
			        8156 => x"00000000",		-- colors: 40, 40, 40, 40
			        8157 => x"00000000",		-- colors: 40, 40, 40, 40
			        8158 => x"00000000",		-- colors: 40, 40, 40, 40
			        8159 => x"00000000",		-- colors: 40, 40, 40, 40
			        8160 => x"00000000",		-- colors: 40, 40, 40, 40
			        8161 => x"00000000",		-- colors: 40, 40, 40, 40
			        8162 => x"00000000",		-- colors: 40, 40, 40, 40
			        8163 => x"00000000",		-- colors: 40, 40, 40, 40
			        8164 => x"00000000",		-- colors: 40, 40, 40, 40
			        8165 => x"00000000",		-- colors: 40, 40, 40, 40
			        8166 => x"00000000",		-- colors: 40, 40, 40, 40
			        8167 => x"00000000",		-- colors: 40, 40, 40, 40
			        8168 => x"00000000",		-- colors: 40, 40, 40, 40
			        8169 => x"00000000",		-- colors: 40, 40, 40, 40
			        8170 => x"00000000",		-- colors: 40, 40, 40, 40
			        8171 => x"00000000",		-- colors: 40, 40, 40, 40
			        8172 => x"00000000",		-- colors: 40, 40, 40, 40
			        8173 => x"00000000",		-- colors: 40, 40, 40, 40
			        8174 => x"00000000",		-- colors: 40, 40, 40, 40
			        8175 => x"00000000",		-- colors: 40, 40, 40, 40
			        8176 => x"00000000",		-- colors: 40, 40, 40, 40
			        8177 => x"00000000",		-- colors: 40, 40, 40, 40
			        8178 => x"00000000",		-- colors: 40, 40, 40, 40
			        8179 => x"00000000",		-- colors: 40, 40, 40, 40
			        8180 => x"00000000",		-- colors: 40, 40, 40, 40
			        8181 => x"00000000",		-- colors: 40, 40, 40, 40
			        8182 => x"00000000",		-- colors: 40, 40, 40, 40
			        8183 => x"00000000",		-- colors: 40, 40, 40, 40
			        8184 => x"00000000",		-- colors: 40, 40, 40, 40
			        8185 => x"00000000",		-- colors: 40, 40, 40, 40
			        8186 => x"00000000",		-- colors: 40, 40, 40, 40
			        8187 => x"00000000",		-- colors: 40, 40, 40, 40
			        8188 => x"00000000",		-- colors: 40, 40, 40, 40
			        8189 => x"00000000",		-- colors: 40, 40, 40, 40
			        8190 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 124
			        8191 => x"00000000",		-- colors: 40, 40, 40, 40
			        8192 => x"00000000",		-- colors: 40, 40, 40, 40
			        8193 => x"00000000",		-- colors: 40, 40, 40, 40
			        8194 => x"00000000",		-- colors: 40, 40, 40, 40
			        8195 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8196 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8197 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8198 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8199 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8200 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8201 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8202 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8203 => x"00000000",		-- colors: 40, 40, 40, 40
			        8204 => x"00000000",		-- colors: 40, 40, 40, 40
			        8205 => x"00000000",		-- colors: 40, 40, 40, 40
			        8206 => x"00000000",		-- colors: 40, 40, 40, 40
			        8207 => x"00000000",		-- colors: 40, 40, 40, 40
			        8208 => x"00000000",		-- colors: 40, 40, 40, 40
			        8209 => x"00000000",		-- colors: 40, 40, 40, 40
			        8210 => x"00000000",		-- colors: 40, 40, 40, 40
			        8211 => x"00000000",		-- colors: 40, 40, 40, 40
			        8212 => x"00000000",		-- colors: 40, 40, 40, 40
			        8213 => x"00000000",		-- colors: 40, 40, 40, 40
			        8214 => x"00000000",		-- colors: 40, 40, 40, 40
			        8215 => x"00000000",		-- colors: 40, 40, 40, 40
			        8216 => x"00000000",		-- colors: 40, 40, 40, 40
			        8217 => x"00000000",		-- colors: 40, 40, 40, 40
			        8218 => x"00000000",		-- colors: 40, 40, 40, 40
			        8219 => x"00000000",		-- colors: 40, 40, 40, 40
			        8220 => x"00000000",		-- colors: 40, 40, 40, 40
			        8221 => x"00000000",		-- colors: 40, 40, 40, 40
			        8222 => x"00000000",		-- colors: 40, 40, 40, 40
			        8223 => x"00000000",		-- colors: 40, 40, 40, 40
			        8224 => x"00000000",		-- colors: 40, 40, 40, 40
			        8225 => x"00000000",		-- colors: 40, 40, 40, 40
			        8226 => x"00000000",		-- colors: 40, 40, 40, 40
			        8227 => x"00000000",		-- colors: 40, 40, 40, 40
			        8228 => x"00000000",		-- colors: 40, 40, 40, 40
			        8229 => x"00000000",		-- colors: 40, 40, 40, 40
			        8230 => x"00000000",		-- colors: 40, 40, 40, 40
			        8231 => x"00000000",		-- colors: 40, 40, 40, 40
			        8232 => x"00000000",		-- colors: 40, 40, 40, 40
			        8233 => x"00000000",		-- colors: 40, 40, 40, 40
			        8234 => x"00000000",		-- colors: 40, 40, 40, 40
			        8235 => x"00000000",		-- colors: 40, 40, 40, 40
			        8236 => x"00000000",		-- colors: 40, 40, 40, 40
			        8237 => x"00000000",		-- colors: 40, 40, 40, 40
			        8238 => x"00000000",		-- colors: 40, 40, 40, 40
			        8239 => x"00000000",		-- colors: 40, 40, 40, 40
			        8240 => x"00000000",		-- colors: 40, 40, 40, 40
			        8241 => x"00000000",		-- colors: 40, 40, 40, 40
			        8242 => x"00000000",		-- colors: 40, 40, 40, 40
			        8243 => x"00000000",		-- colors: 40, 40, 40, 40
			        8244 => x"00000000",		-- colors: 40, 40, 40, 40
			        8245 => x"00000000",		-- colors: 40, 40, 40, 40
			        8246 => x"00000000",		-- colors: 40, 40, 40, 40
			        8247 => x"00000000",		-- colors: 40, 40, 40, 40
			        8248 => x"00000000",		-- colors: 40, 40, 40, 40
			        8249 => x"00000000",		-- colors: 40, 40, 40, 40
			        8250 => x"00000000",		-- colors: 40, 40, 40, 40
			        8251 => x"00000000",		-- colors: 40, 40, 40, 40
			        8252 => x"00000000",		-- colors: 40, 40, 40, 40
			        8253 => x"00000000",		-- colors: 40, 40, 40, 40
			        8254 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 125
			        8255 => x"00000000",		-- colors: 40, 40, 40, 40
			        8256 => x"00000000",		-- colors: 40, 40, 40, 40
			        8257 => x"00000000",		-- colors: 40, 40, 40, 40
			        8258 => x"00000000",		-- colors: 40, 40, 40, 40
			        8259 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8260 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8261 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8262 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8263 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8264 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8265 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8266 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8267 => x"00000000",		-- colors: 40, 40, 40, 40
			        8268 => x"00000000",		-- colors: 40, 40, 40, 40
			        8269 => x"00000000",		-- colors: 40, 40, 40, 40
			        8270 => x"00000000",		-- colors: 40, 40, 40, 40
			        8271 => x"00000000",		-- colors: 40, 40, 40, 40
			        8272 => x"00000000",		-- colors: 40, 40, 40, 40
			        8273 => x"00000000",		-- colors: 40, 40, 40, 40
			        8274 => x"00000000",		-- colors: 40, 40, 40, 40
			        8275 => x"00000000",		-- colors: 40, 40, 40, 40
			        8276 => x"00000000",		-- colors: 40, 40, 40, 40
			        8277 => x"00000000",		-- colors: 40, 40, 40, 40
			        8278 => x"00000000",		-- colors: 40, 40, 40, 40
			        8279 => x"00000000",		-- colors: 40, 40, 40, 40
			        8280 => x"00000000",		-- colors: 40, 40, 40, 40
			        8281 => x"00000000",		-- colors: 40, 40, 40, 40
			        8282 => x"00000000",		-- colors: 40, 40, 40, 40
			        8283 => x"00000000",		-- colors: 40, 40, 40, 40
			        8284 => x"00000000",		-- colors: 40, 40, 40, 40
			        8285 => x"00000000",		-- colors: 40, 40, 40, 40
			        8286 => x"00000000",		-- colors: 40, 40, 40, 40
			        8287 => x"00000000",		-- colors: 40, 40, 40, 40
			        8288 => x"00000000",		-- colors: 40, 40, 40, 40
			        8289 => x"00000000",		-- colors: 40, 40, 40, 40
			        8290 => x"00000000",		-- colors: 40, 40, 40, 40
			        8291 => x"00000000",		-- colors: 40, 40, 40, 40
			        8292 => x"00000000",		-- colors: 40, 40, 40, 40
			        8293 => x"00000000",		-- colors: 40, 40, 40, 40
			        8294 => x"00000000",		-- colors: 40, 40, 40, 40
			        8295 => x"00000000",		-- colors: 40, 40, 40, 40
			        8296 => x"00000000",		-- colors: 40, 40, 40, 40
			        8297 => x"00000000",		-- colors: 40, 40, 40, 40
			        8298 => x"00000000",		-- colors: 40, 40, 40, 40
			        8299 => x"00000000",		-- colors: 40, 40, 40, 40
			        8300 => x"00000000",		-- colors: 40, 40, 40, 40
			        8301 => x"00000000",		-- colors: 40, 40, 40, 40
			        8302 => x"00000000",		-- colors: 40, 40, 40, 40
			        8303 => x"00000000",		-- colors: 40, 40, 40, 40
			        8304 => x"00000000",		-- colors: 40, 40, 40, 40
			        8305 => x"00000000",		-- colors: 40, 40, 40, 40
			        8306 => x"00000000",		-- colors: 40, 40, 40, 40
			        8307 => x"00000000",		-- colors: 40, 40, 40, 40
			        8308 => x"00000000",		-- colors: 40, 40, 40, 40
			        8309 => x"00000000",		-- colors: 40, 40, 40, 40
			        8310 => x"00000000",		-- colors: 40, 40, 40, 40
			        8311 => x"00000000",		-- colors: 40, 40, 40, 40
			        8312 => x"00000000",		-- colors: 40, 40, 40, 40
			        8313 => x"00000000",		-- colors: 40, 40, 40, 40
			        8314 => x"00000000",		-- colors: 40, 40, 40, 40
			        8315 => x"00000000",		-- colors: 40, 40, 40, 40
			        8316 => x"00000000",		-- colors: 40, 40, 40, 40
			        8317 => x"00000000",		-- colors: 40, 40, 40, 40
			        8318 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 126
			        8319 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8320 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8321 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8322 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8323 => x"00000000",		-- colors: 40, 40, 40, 40
			        8324 => x"00000000",		-- colors: 40, 40, 40, 40
			        8325 => x"00000000",		-- colors: 40, 40, 40, 40
			        8326 => x"00000000",		-- colors: 40, 40, 40, 40
			        8327 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8328 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8329 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8330 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8331 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8332 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8333 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8334 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8335 => x"00000000",		-- colors: 40, 40, 40, 40
			        8336 => x"00000000",		-- colors: 40, 40, 40, 40
			        8337 => x"00000000",		-- colors: 40, 40, 40, 40
			        8338 => x"00000000",		-- colors: 40, 40, 40, 40
			        8339 => x"00000000",		-- colors: 40, 40, 40, 40
			        8340 => x"00000000",		-- colors: 40, 40, 40, 40
			        8341 => x"00000000",		-- colors: 40, 40, 40, 40
			        8342 => x"00000000",		-- colors: 40, 40, 40, 40
			        8343 => x"00000000",		-- colors: 40, 40, 40, 40
			        8344 => x"00000000",		-- colors: 40, 40, 40, 40
			        8345 => x"00000000",		-- colors: 40, 40, 40, 40
			        8346 => x"00000000",		-- colors: 40, 40, 40, 40
			        8347 => x"00000000",		-- colors: 40, 40, 40, 40
			        8348 => x"00000000",		-- colors: 40, 40, 40, 40
			        8349 => x"00000000",		-- colors: 40, 40, 40, 40
			        8350 => x"00000000",		-- colors: 40, 40, 40, 40
			        8351 => x"00000000",		-- colors: 40, 40, 40, 40
			        8352 => x"00000000",		-- colors: 40, 40, 40, 40
			        8353 => x"00000000",		-- colors: 40, 40, 40, 40
			        8354 => x"00000000",		-- colors: 40, 40, 40, 40
			        8355 => x"00000000",		-- colors: 40, 40, 40, 40
			        8356 => x"00000000",		-- colors: 40, 40, 40, 40
			        8357 => x"00000000",		-- colors: 40, 40, 40, 40
			        8358 => x"00000000",		-- colors: 40, 40, 40, 40
			        8359 => x"00000000",		-- colors: 40, 40, 40, 40
			        8360 => x"00000000",		-- colors: 40, 40, 40, 40
			        8361 => x"00000000",		-- colors: 40, 40, 40, 40
			        8362 => x"00000000",		-- colors: 40, 40, 40, 40
			        8363 => x"00000000",		-- colors: 40, 40, 40, 40
			        8364 => x"00000000",		-- colors: 40, 40, 40, 40
			        8365 => x"00000000",		-- colors: 40, 40, 40, 40
			        8366 => x"00000000",		-- colors: 40, 40, 40, 40
			        8367 => x"00000000",		-- colors: 40, 40, 40, 40
			        8368 => x"00000000",		-- colors: 40, 40, 40, 40
			        8369 => x"00000000",		-- colors: 40, 40, 40, 40
			        8370 => x"00000000",		-- colors: 40, 40, 40, 40
			        8371 => x"00000000",		-- colors: 40, 40, 40, 40
			        8372 => x"00000000",		-- colors: 40, 40, 40, 40
			        8373 => x"00000000",		-- colors: 40, 40, 40, 40
			        8374 => x"00000000",		-- colors: 40, 40, 40, 40
			        8375 => x"00000000",		-- colors: 40, 40, 40, 40
			        8376 => x"00000000",		-- colors: 40, 40, 40, 40
			        8377 => x"00000000",		-- colors: 40, 40, 40, 40
			        8378 => x"00000000",		-- colors: 40, 40, 40, 40
			        8379 => x"00000000",		-- colors: 40, 40, 40, 40
			        8380 => x"00000000",		-- colors: 40, 40, 40, 40
			        8381 => x"00000000",		-- colors: 40, 40, 40, 40
			        8382 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 127
			        8383 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8384 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8385 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8386 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8387 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8388 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8389 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8390 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8391 => x"00000000",		-- colors: 40, 40, 40, 40
			        8392 => x"00000000",		-- colors: 40, 40, 40, 40
			        8393 => x"00000000",		-- colors: 40, 40, 40, 40
			        8394 => x"00000000",		-- colors: 40, 40, 40, 40
			        8395 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8396 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8397 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8398 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8399 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8400 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8401 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8402 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8403 => x"00000000",		-- colors: 40, 40, 40, 40
			        8404 => x"00000000",		-- colors: 40, 40, 40, 40
			        8405 => x"00000000",		-- colors: 40, 40, 40, 40
			        8406 => x"00000000",		-- colors: 40, 40, 40, 40
			        8407 => x"32323232",		-- colors: 50, 50, 50, 50
			        8408 => x"32323232",		-- colors: 50, 50, 50, 50
			        8409 => x"32323232",		-- colors: 50, 50, 50, 50
			        8410 => x"32323232",		-- colors: 50, 50, 50, 50
			        8411 => x"00000000",		-- colors: 40, 40, 40, 40
			        8412 => x"00000000",		-- colors: 40, 40, 40, 40
			        8413 => x"00000000",		-- colors: 40, 40, 40, 40
			        8414 => x"00000000",		-- colors: 40, 40, 40, 40
			        8415 => x"00000000",		-- colors: 40, 40, 40, 40
			        8416 => x"00000000",		-- colors: 40, 40, 40, 40
			        8417 => x"00000000",		-- colors: 40, 40, 40, 40
			        8418 => x"00000000",		-- colors: 40, 40, 40, 40
			        8419 => x"00000000",		-- colors: 40, 40, 40, 40
			        8420 => x"00000000",		-- colors: 40, 40, 40, 40
			        8421 => x"00000000",		-- colors: 40, 40, 40, 40
			        8422 => x"00000000",		-- colors: 40, 40, 40, 40
			        8423 => x"32323232",		-- colors: 50, 50, 50, 50
			        8424 => x"32323232",		-- colors: 50, 50, 50, 50
			        8425 => x"32323232",		-- colors: 50, 50, 50, 50
			        8426 => x"32323232",		-- colors: 50, 50, 50, 50
			        8427 => x"00000000",		-- colors: 40, 40, 40, 40
			        8428 => x"00000000",		-- colors: 40, 40, 40, 40
			        8429 => x"00000000",		-- colors: 40, 40, 40, 40
			        8430 => x"00000000",		-- colors: 40, 40, 40, 40
			        8431 => x"00000000",		-- colors: 40, 40, 40, 40
			        8432 => x"00000000",		-- colors: 40, 40, 40, 40
			        8433 => x"00000000",		-- colors: 40, 40, 40, 40
			        8434 => x"00000000",		-- colors: 40, 40, 40, 40
			        8435 => x"00000000",		-- colors: 40, 40, 40, 40
			        8436 => x"00000000",		-- colors: 40, 40, 40, 40
			        8437 => x"00000000",		-- colors: 40, 40, 40, 40
			        8438 => x"00000000",		-- colors: 40, 40, 40, 40
			        8439 => x"32323232",		-- colors: 50, 50, 50, 50
			        8440 => x"32323232",		-- colors: 50, 50, 50, 50
			        8441 => x"32323232",		-- colors: 50, 50, 50, 50
			        8442 => x"32323232",		-- colors: 50, 50, 50, 50
			        8443 => x"00000000",		-- colors: 40, 40, 40, 40
			        8444 => x"00000000",		-- colors: 40, 40, 40, 40
			        8445 => x"00000000",		-- colors: 40, 40, 40, 40
			        8446 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 128
			        8447 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8448 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8449 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8450 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8451 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8452 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8453 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8454 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8455 => x"00000000",		-- colors: 40, 40, 40, 40
			        8456 => x"00000000",		-- colors: 40, 40, 40, 40
			        8457 => x"00000000",		-- colors: 40, 40, 40, 40
			        8458 => x"00000000",		-- colors: 40, 40, 40, 40
			        8459 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8460 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8461 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8462 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8463 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8464 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8465 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8466 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8467 => x"00000000",		-- colors: 40, 40, 40, 40
			        8468 => x"00000000",		-- colors: 40, 40, 40, 40
			        8469 => x"00000000",		-- colors: 40, 40, 40, 40
			        8470 => x"00000000",		-- colors: 40, 40, 40, 40
			        8471 => x"00000000",		-- colors: 40, 40, 40, 40
			        8472 => x"00000000",		-- colors: 40, 40, 40, 40
			        8473 => x"00000000",		-- colors: 40, 40, 40, 40
			        8474 => x"00000000",		-- colors: 40, 40, 40, 40
			        8475 => x"00000000",		-- colors: 40, 40, 40, 40
			        8476 => x"00000000",		-- colors: 40, 40, 40, 40
			        8477 => x"00000000",		-- colors: 40, 40, 40, 40
			        8478 => x"00000000",		-- colors: 40, 40, 40, 40
			        8479 => x"00000000",		-- colors: 40, 40, 40, 40
			        8480 => x"00000000",		-- colors: 40, 40, 40, 40
			        8481 => x"00000000",		-- colors: 40, 40, 40, 40
			        8482 => x"00000000",		-- colors: 40, 40, 40, 40
			        8483 => x"00000000",		-- colors: 40, 40, 40, 40
			        8484 => x"00000000",		-- colors: 40, 40, 40, 40
			        8485 => x"00000000",		-- colors: 40, 40, 40, 40
			        8486 => x"00000000",		-- colors: 40, 40, 40, 40
			        8487 => x"00000000",		-- colors: 40, 40, 40, 40
			        8488 => x"00000000",		-- colors: 40, 40, 40, 40
			        8489 => x"00000000",		-- colors: 40, 40, 40, 40
			        8490 => x"00000000",		-- colors: 40, 40, 40, 40
			        8491 => x"00000000",		-- colors: 40, 40, 40, 40
			        8492 => x"00000000",		-- colors: 40, 40, 40, 40
			        8493 => x"00000000",		-- colors: 40, 40, 40, 40
			        8494 => x"00000000",		-- colors: 40, 40, 40, 40
			        8495 => x"00000000",		-- colors: 40, 40, 40, 40
			        8496 => x"00000000",		-- colors: 40, 40, 40, 40
			        8497 => x"00000000",		-- colors: 40, 40, 40, 40
			        8498 => x"00000000",		-- colors: 40, 40, 40, 40
			        8499 => x"00000000",		-- colors: 40, 40, 40, 40
			        8500 => x"00000000",		-- colors: 40, 40, 40, 40
			        8501 => x"00000000",		-- colors: 40, 40, 40, 40
			        8502 => x"00000000",		-- colors: 40, 40, 40, 40
			        8503 => x"00000000",		-- colors: 40, 40, 40, 40
			        8504 => x"00000000",		-- colors: 40, 40, 40, 40
			        8505 => x"00000000",		-- colors: 40, 40, 40, 40
			        8506 => x"00000000",		-- colors: 40, 40, 40, 40
			        8507 => x"00000000",		-- colors: 40, 40, 40, 40
			        8508 => x"00000000",		-- colors: 40, 40, 40, 40
			        8509 => x"00000000",		-- colors: 40, 40, 40, 40
			        8510 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 129
			        8511 => x"00000000",		-- colors: 40, 40, 40, 40
			        8512 => x"00000000",		-- colors: 40, 40, 40, 40
			        8513 => x"00000000",		-- colors: 40, 40, 40, 40
			        8514 => x"00000000",		-- colors: 40, 40, 40, 40
			        8515 => x"00000000",		-- colors: 40, 40, 40, 40
			        8516 => x"00000000",		-- colors: 40, 40, 40, 40
			        8517 => x"00000000",		-- colors: 40, 40, 40, 40
			        8518 => x"00000000",		-- colors: 40, 40, 40, 40
			        8519 => x"00000000",		-- colors: 40, 40, 40, 40
			        8520 => x"00000000",		-- colors: 40, 40, 40, 40
			        8521 => x"00000000",		-- colors: 40, 40, 40, 40
			        8522 => x"00000000",		-- colors: 40, 40, 40, 40
			        8523 => x"00000000",		-- colors: 40, 40, 40, 40
			        8524 => x"00000000",		-- colors: 40, 40, 40, 40
			        8525 => x"00000000",		-- colors: 40, 40, 40, 40
			        8526 => x"00000000",		-- colors: 40, 40, 40, 40
			        8527 => x"00000000",		-- colors: 40, 40, 40, 40
			        8528 => x"00000000",		-- colors: 40, 40, 40, 40
			        8529 => x"00000000",		-- colors: 40, 40, 40, 40
			        8530 => x"00000000",		-- colors: 40, 40, 40, 40
			        8531 => x"00000000",		-- colors: 40, 40, 40, 40
			        8532 => x"00000000",		-- colors: 40, 40, 40, 40
			        8533 => x"00000000",		-- colors: 40, 40, 40, 40
			        8534 => x"00000000",		-- colors: 40, 40, 40, 40
			        8535 => x"00000000",		-- colors: 40, 40, 40, 40
			        8536 => x"00000000",		-- colors: 40, 40, 40, 40
			        8537 => x"00000000",		-- colors: 40, 40, 40, 40
			        8538 => x"00000000",		-- colors: 40, 40, 40, 40
			        8539 => x"00000000",		-- colors: 40, 40, 40, 40
			        8540 => x"00000000",		-- colors: 40, 40, 40, 40
			        8541 => x"00000000",		-- colors: 40, 40, 40, 40
			        8542 => x"00000000",		-- colors: 40, 40, 40, 40
			        8543 => x"00000000",		-- colors: 40, 40, 40, 40
			        8544 => x"00000000",		-- colors: 40, 40, 40, 40
			        8545 => x"00000000",		-- colors: 40, 40, 40, 40
			        8546 => x"00000000",		-- colors: 40, 40, 40, 40
			        8547 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8548 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8549 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8550 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8551 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8552 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8553 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8554 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8555 => x"00000000",		-- colors: 40, 40, 40, 40
			        8556 => x"00000000",		-- colors: 40, 40, 40, 40
			        8557 => x"00000000",		-- colors: 40, 40, 40, 40
			        8558 => x"00000000",		-- colors: 40, 40, 40, 40
			        8559 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8560 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8561 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8562 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8563 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8564 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8565 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8566 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8567 => x"00000000",		-- colors: 40, 40, 40, 40
			        8568 => x"00000000",		-- colors: 40, 40, 40, 40
			        8569 => x"00000000",		-- colors: 40, 40, 40, 40
			        8570 => x"00000000",		-- colors: 40, 40, 40, 40
			        8571 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8572 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8573 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8574 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60

			                --  sprite 130
			        8575 => x"00000000",		-- colors: 40, 40, 40, 40
			        8576 => x"00000000",		-- colors: 40, 40, 40, 40
			        8577 => x"00000000",		-- colors: 40, 40, 40, 40
			        8578 => x"00000000",		-- colors: 40, 40, 40, 40
			        8579 => x"00000000",		-- colors: 40, 40, 40, 40
			        8580 => x"00000000",		-- colors: 40, 40, 40, 40
			        8581 => x"00000000",		-- colors: 40, 40, 40, 40
			        8582 => x"00000000",		-- colors: 40, 40, 40, 40
			        8583 => x"00000000",		-- colors: 40, 40, 40, 40
			        8584 => x"00000000",		-- colors: 40, 40, 40, 40
			        8585 => x"00000000",		-- colors: 40, 40, 40, 40
			        8586 => x"00000000",		-- colors: 40, 40, 40, 40
			        8587 => x"00000000",		-- colors: 40, 40, 40, 40
			        8588 => x"00000000",		-- colors: 40, 40, 40, 40
			        8589 => x"00000000",		-- colors: 40, 40, 40, 40
			        8590 => x"00000000",		-- colors: 40, 40, 40, 40
			        8591 => x"00000000",		-- colors: 40, 40, 40, 40
			        8592 => x"00000000",		-- colors: 40, 40, 40, 40
			        8593 => x"00000000",		-- colors: 40, 40, 40, 40
			        8594 => x"00000000",		-- colors: 40, 40, 40, 40
			        8595 => x"00000000",		-- colors: 40, 40, 40, 40
			        8596 => x"00000000",		-- colors: 40, 40, 40, 40
			        8597 => x"00000000",		-- colors: 40, 40, 40, 40
			        8598 => x"00000000",		-- colors: 40, 40, 40, 40
			        8599 => x"00000000",		-- colors: 40, 40, 40, 40
			        8600 => x"00000000",		-- colors: 40, 40, 40, 40
			        8601 => x"00000000",		-- colors: 40, 40, 40, 40
			        8602 => x"00000000",		-- colors: 40, 40, 40, 40
			        8603 => x"00000000",		-- colors: 40, 40, 40, 40
			        8604 => x"00000000",		-- colors: 40, 40, 40, 40
			        8605 => x"00000000",		-- colors: 40, 40, 40, 40
			        8606 => x"00000000",		-- colors: 40, 40, 40, 40
			        8607 => x"00000000",		-- colors: 40, 40, 40, 40
			        8608 => x"00000000",		-- colors: 40, 40, 40, 40
			        8609 => x"00000000",		-- colors: 40, 40, 40, 40
			        8610 => x"00000000",		-- colors: 40, 40, 40, 40
			        8611 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8612 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8613 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8614 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8615 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8616 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8617 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8618 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8619 => x"00000000",		-- colors: 40, 40, 40, 40
			        8620 => x"00000000",		-- colors: 40, 40, 40, 40
			        8621 => x"00000000",		-- colors: 40, 40, 40, 40
			        8622 => x"00000000",		-- colors: 40, 40, 40, 40
			        8623 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8624 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8625 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8626 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8627 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8628 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8629 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8630 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8631 => x"00000000",		-- colors: 40, 40, 40, 40
			        8632 => x"00000000",		-- colors: 40, 40, 40, 40
			        8633 => x"00000000",		-- colors: 40, 40, 40, 40
			        8634 => x"00000000",		-- colors: 40, 40, 40, 40
			        8635 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8636 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8637 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8638 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60

			                --  sprite 131
			        8639 => x"32323232",		-- colors: 50, 50, 50, 50
			        8640 => x"32323232",		-- colors: 50, 50, 50, 50
			        8641 => x"32323232",		-- colors: 50, 50, 50, 50
			        8642 => x"32323232",		-- colors: 50, 50, 50, 50
			        8643 => x"32323232",		-- colors: 50, 50, 50, 50
			        8644 => x"32323232",		-- colors: 50, 50, 50, 50
			        8645 => x"32323232",		-- colors: 50, 50, 50, 50
			        8646 => x"32323232",		-- colors: 50, 50, 50, 50
			        8647 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
			        8648 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
			        8649 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
			        8650 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
			        8651 => x"32323232",		-- colors: 50, 50, 50, 50
			        8652 => x"32323232",		-- colors: 50, 50, 50, 50
			        8653 => x"32323232",		-- colors: 50, 50, 50, 50
			        8654 => x"32323232",		-- colors: 50, 50, 50, 50
			        8655 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
			        8656 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
			        8657 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
			        8658 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
			        8659 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
			        8660 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
			        8661 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
			        8662 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
			        8663 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
			        8664 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
			        8665 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
			        8666 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
			        8667 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
			        8668 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
			        8669 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
			        8670 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
			        8671 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
			        8672 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
			        8673 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
			        8674 => x"3E3E3E3E",		-- colors: 62, 62, 62, 62
			        8675 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8676 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8677 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8678 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8679 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8680 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8681 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8682 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8683 => x"00000000",		-- colors: 40, 40, 40, 40
			        8684 => x"00000000",		-- colors: 40, 40, 40, 40
			        8685 => x"00000000",		-- colors: 40, 40, 40, 40
			        8686 => x"00000000",		-- colors: 40, 40, 40, 40
			        8687 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8688 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8689 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8690 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8691 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8692 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8693 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8694 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8695 => x"00000000",		-- colors: 40, 40, 40, 40
			        8696 => x"00000000",		-- colors: 40, 40, 40, 40
			        8697 => x"00000000",		-- colors: 40, 40, 40, 40
			        8698 => x"00000000",		-- colors: 40, 40, 40, 40
			        8699 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8700 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8701 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8702 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60

			                --  sprite 132
			        8703 => x"00000000",		-- colors: 40, 40, 40, 40
			        8704 => x"00000000",		-- colors: 40, 40, 40, 40
			        8705 => x"00000000",		-- colors: 40, 40, 40, 40
			        8706 => x"00000000",		-- colors: 40, 40, 40, 40
			        8707 => x"00000000",		-- colors: 40, 40, 40, 40
			        8708 => x"00000000",		-- colors: 40, 40, 40, 40
			        8709 => x"00000000",		-- colors: 40, 40, 40, 40
			        8710 => x"00000000",		-- colors: 40, 40, 40, 40
			        8711 => x"00000000",		-- colors: 40, 40, 40, 40
			        8712 => x"00000000",		-- colors: 40, 40, 40, 40
			        8713 => x"00000000",		-- colors: 40, 40, 40, 40
			        8714 => x"00000000",		-- colors: 40, 40, 40, 40
			        8715 => x"00000000",		-- colors: 40, 40, 40, 40
			        8716 => x"00000000",		-- colors: 40, 40, 40, 40
			        8717 => x"00000000",		-- colors: 40, 40, 40, 40
			        8718 => x"00000000",		-- colors: 40, 40, 40, 40
			        8719 => x"00000000",		-- colors: 40, 40, 40, 40
			        8720 => x"00000000",		-- colors: 40, 40, 40, 40
			        8721 => x"00000000",		-- colors: 40, 40, 40, 40
			        8722 => x"00000000",		-- colors: 40, 40, 40, 40
			        8723 => x"00000000",		-- colors: 40, 40, 40, 40
			        8724 => x"00000000",		-- colors: 40, 40, 40, 40
			        8725 => x"00000000",		-- colors: 40, 40, 40, 40
			        8726 => x"00000000",		-- colors: 40, 40, 40, 40
			        8727 => x"00000000",		-- colors: 40, 40, 40, 40
			        8728 => x"00000000",		-- colors: 40, 40, 40, 40
			        8729 => x"00000000",		-- colors: 40, 40, 40, 40
			        8730 => x"00000000",		-- colors: 40, 40, 40, 40
			        8731 => x"00000000",		-- colors: 40, 40, 40, 40
			        8732 => x"00000000",		-- colors: 40, 40, 40, 40
			        8733 => x"00000000",		-- colors: 40, 40, 40, 40
			        8734 => x"00000000",		-- colors: 40, 40, 40, 40
			        8735 => x"00000000",		-- colors: 40, 40, 40, 40
			        8736 => x"00000000",		-- colors: 40, 40, 40, 40
			        8737 => x"00000000",		-- colors: 40, 40, 40, 40
			        8738 => x"00000000",		-- colors: 40, 40, 40, 40
			        8739 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8740 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8741 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8742 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8743 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8744 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8745 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8746 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8747 => x"00000000",		-- colors: 40, 40, 40, 40
			        8748 => x"00000000",		-- colors: 40, 40, 40, 40
			        8749 => x"00000000",		-- colors: 40, 40, 40, 40
			        8750 => x"00000000",		-- colors: 40, 40, 40, 40
			        8751 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8752 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8753 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8754 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8755 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8756 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8757 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8758 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8759 => x"00000000",		-- colors: 40, 40, 40, 40
			        8760 => x"00000000",		-- colors: 40, 40, 40, 40
			        8761 => x"00000000",		-- colors: 40, 40, 40, 40
			        8762 => x"00000000",		-- colors: 40, 40, 40, 40
			        8763 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8764 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8765 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8766 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60

			                --  sprite 133
			        8767 => x"00000000",		-- colors: 40, 40, 40, 40
			        8768 => x"00000000",		-- colors: 40, 40, 40, 40
			        8769 => x"00000000",		-- colors: 40, 40, 40, 40
			        8770 => x"00000000",		-- colors: 40, 40, 40, 40
			        8771 => x"00000000",		-- colors: 40, 40, 40, 40
			        8772 => x"00000000",		-- colors: 40, 40, 40, 40
			        8773 => x"00000000",		-- colors: 40, 40, 40, 40
			        8774 => x"00000000",		-- colors: 40, 40, 40, 40
			        8775 => x"00000000",		-- colors: 40, 40, 40, 40
			        8776 => x"00000000",		-- colors: 40, 40, 40, 40
			        8777 => x"00000000",		-- colors: 40, 40, 40, 40
			        8778 => x"00000000",		-- colors: 40, 40, 40, 40
			        8779 => x"00000000",		-- colors: 40, 40, 40, 40
			        8780 => x"00000000",		-- colors: 40, 40, 40, 40
			        8781 => x"00000000",		-- colors: 40, 40, 40, 40
			        8782 => x"00000000",		-- colors: 40, 40, 40, 40
			        8783 => x"00000000",		-- colors: 40, 40, 40, 40
			        8784 => x"00000000",		-- colors: 40, 40, 40, 40
			        8785 => x"00000000",		-- colors: 40, 40, 40, 40
			        8786 => x"00000000",		-- colors: 40, 40, 40, 40
			        8787 => x"00000000",		-- colors: 40, 40, 40, 40
			        8788 => x"00000000",		-- colors: 40, 40, 40, 40
			        8789 => x"00000000",		-- colors: 40, 40, 40, 40
			        8790 => x"00000000",		-- colors: 40, 40, 40, 40
			        8791 => x"00000000",		-- colors: 40, 40, 40, 40
			        8792 => x"00000000",		-- colors: 40, 40, 40, 40
			        8793 => x"00000000",		-- colors: 40, 40, 40, 40
			        8794 => x"00000000",		-- colors: 40, 40, 40, 40
			        8795 => x"00000000",		-- colors: 40, 40, 40, 40
			        8796 => x"00000000",		-- colors: 40, 40, 40, 40
			        8797 => x"00000000",		-- colors: 40, 40, 40, 40
			        8798 => x"00000000",		-- colors: 40, 40, 40, 40
			        8799 => x"00000000",		-- colors: 40, 40, 40, 40
			        8800 => x"00000000",		-- colors: 40, 40, 40, 40
			        8801 => x"00000000",		-- colors: 40, 40, 40, 40
			        8802 => x"00000000",		-- colors: 40, 40, 40, 40
			        8803 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8804 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8805 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8806 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8807 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8808 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8809 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8810 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8811 => x"00000000",		-- colors: 40, 40, 40, 40
			        8812 => x"00000000",		-- colors: 40, 40, 40, 40
			        8813 => x"00000000",		-- colors: 40, 40, 40, 40
			        8814 => x"00000000",		-- colors: 40, 40, 40, 40
			        8815 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8816 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8817 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8818 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8819 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8820 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8821 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8822 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8823 => x"00000000",		-- colors: 40, 40, 40, 40
			        8824 => x"00000000",		-- colors: 40, 40, 40, 40
			        8825 => x"00000000",		-- colors: 40, 40, 40, 40
			        8826 => x"00000000",		-- colors: 40, 40, 40, 40
			        8827 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8828 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8829 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8830 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60

			                --  sprite 134
			        8831 => x"00000000",		-- colors: 40, 40, 40, 40
			        8832 => x"00000000",		-- colors: 40, 40, 40, 40
			        8833 => x"00000000",		-- colors: 40, 40, 40, 40
			        8834 => x"00000000",		-- colors: 40, 40, 40, 40
			        8835 => x"00000000",		-- colors: 40, 40, 40, 40
			        8836 => x"00000000",		-- colors: 40, 40, 40, 40
			        8837 => x"00000000",		-- colors: 40, 40, 40, 40
			        8838 => x"00000000",		-- colors: 40, 40, 40, 40
			        8839 => x"00000000",		-- colors: 40, 40, 40, 40
			        8840 => x"00000000",		-- colors: 40, 40, 40, 40
			        8841 => x"00000000",		-- colors: 40, 40, 40, 40
			        8842 => x"00000000",		-- colors: 40, 40, 40, 40
			        8843 => x"00000000",		-- colors: 40, 40, 40, 40
			        8844 => x"00000000",		-- colors: 40, 40, 40, 40
			        8845 => x"00000000",		-- colors: 40, 40, 40, 40
			        8846 => x"00000000",		-- colors: 40, 40, 40, 40
			        8847 => x"00000000",		-- colors: 40, 40, 40, 40
			        8848 => x"00000000",		-- colors: 40, 40, 40, 40
			        8849 => x"00000000",		-- colors: 40, 40, 40, 40
			        8850 => x"00000000",		-- colors: 40, 40, 40, 40
			        8851 => x"00000000",		-- colors: 40, 40, 40, 40
			        8852 => x"00000000",		-- colors: 40, 40, 40, 40
			        8853 => x"00000000",		-- colors: 40, 40, 40, 40
			        8854 => x"00000000",		-- colors: 40, 40, 40, 40
			        8855 => x"00000000",		-- colors: 40, 40, 40, 40
			        8856 => x"00000000",		-- colors: 40, 40, 40, 40
			        8857 => x"00000000",		-- colors: 40, 40, 40, 40
			        8858 => x"00000000",		-- colors: 40, 40, 40, 40
			        8859 => x"00000000",		-- colors: 40, 40, 40, 40
			        8860 => x"00000000",		-- colors: 40, 40, 40, 40
			        8861 => x"00000000",		-- colors: 40, 40, 40, 40
			        8862 => x"00000000",		-- colors: 40, 40, 40, 40
			        8863 => x"00000000",		-- colors: 40, 40, 40, 40
			        8864 => x"00000000",		-- colors: 40, 40, 40, 40
			        8865 => x"00000000",		-- colors: 40, 40, 40, 40
			        8866 => x"00000000",		-- colors: 40, 40, 40, 40
			        8867 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8868 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8869 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8870 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8871 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8872 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8873 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8874 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8875 => x"00000000",		-- colors: 40, 40, 40, 40
			        8876 => x"00000000",		-- colors: 40, 40, 40, 40
			        8877 => x"00000000",		-- colors: 40, 40, 40, 40
			        8878 => x"00000000",		-- colors: 40, 40, 40, 40
			        8879 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8880 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8881 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8882 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8883 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8884 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8885 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8886 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8887 => x"00000000",		-- colors: 40, 40, 40, 40
			        8888 => x"00000000",		-- colors: 40, 40, 40, 40
			        8889 => x"00000000",		-- colors: 40, 40, 40, 40
			        8890 => x"00000000",		-- colors: 40, 40, 40, 40
			        8891 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8892 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8893 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8894 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60

			                --  sprite 135
			        8895 => x"00000000",		-- colors: 40, 40, 40, 40
			        8896 => x"00000000",		-- colors: 40, 40, 40, 40
			        8897 => x"00000000",		-- colors: 40, 40, 40, 40
			        8898 => x"00000000",		-- colors: 40, 40, 40, 40
			        8899 => x"00000000",		-- colors: 40, 40, 40, 40
			        8900 => x"00000000",		-- colors: 40, 40, 40, 40
			        8901 => x"00000000",		-- colors: 40, 40, 40, 40
			        8902 => x"00000000",		-- colors: 40, 40, 40, 40
			        8903 => x"00000000",		-- colors: 40, 40, 40, 40
			        8904 => x"00000000",		-- colors: 40, 40, 40, 40
			        8905 => x"00000000",		-- colors: 40, 40, 40, 40
			        8906 => x"00000000",		-- colors: 40, 40, 40, 40
			        8907 => x"00000000",		-- colors: 40, 40, 40, 40
			        8908 => x"00000000",		-- colors: 40, 40, 40, 40
			        8909 => x"00000000",		-- colors: 40, 40, 40, 40
			        8910 => x"00000000",		-- colors: 40, 40, 40, 40
			        8911 => x"00000000",		-- colors: 40, 40, 40, 40
			        8912 => x"00000000",		-- colors: 40, 40, 40, 40
			        8913 => x"00000000",		-- colors: 40, 40, 40, 40
			        8914 => x"00000000",		-- colors: 40, 40, 40, 40
			        8915 => x"00000000",		-- colors: 40, 40, 40, 40
			        8916 => x"00000000",		-- colors: 40, 40, 40, 40
			        8917 => x"00000000",		-- colors: 40, 40, 40, 40
			        8918 => x"00000000",		-- colors: 40, 40, 40, 40
			        8919 => x"00000000",		-- colors: 40, 40, 40, 40
			        8920 => x"00000000",		-- colors: 40, 40, 40, 40
			        8921 => x"00000000",		-- colors: 40, 40, 40, 40
			        8922 => x"00000000",		-- colors: 40, 40, 40, 40
			        8923 => x"00000000",		-- colors: 40, 40, 40, 40
			        8924 => x"00000000",		-- colors: 40, 40, 40, 40
			        8925 => x"00000000",		-- colors: 40, 40, 40, 40
			        8926 => x"00000000",		-- colors: 40, 40, 40, 40
			        8927 => x"00000000",		-- colors: 40, 40, 40, 40
			        8928 => x"00000000",		-- colors: 40, 40, 40, 40
			        8929 => x"00000000",		-- colors: 40, 40, 40, 40
			        8930 => x"00000000",		-- colors: 40, 40, 40, 40
			        8931 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8932 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8933 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8934 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8935 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8936 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8937 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8938 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8939 => x"00000000",		-- colors: 40, 40, 40, 40
			        8940 => x"00000000",		-- colors: 40, 40, 40, 40
			        8941 => x"00000000",		-- colors: 40, 40, 40, 40
			        8942 => x"00000000",		-- colors: 40, 40, 40, 40
			        8943 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8944 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8945 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8946 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8947 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8948 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8949 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8950 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8951 => x"00000000",		-- colors: 40, 40, 40, 40
			        8952 => x"00000000",		-- colors: 40, 40, 40, 40
			        8953 => x"00000000",		-- colors: 40, 40, 40, 40
			        8954 => x"00000000",		-- colors: 40, 40, 40, 40
			        8955 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8956 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8957 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8958 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60

			                --  sprite 136
			        8959 => x"00000000",		-- colors: 40, 40, 40, 40
			        8960 => x"00000000",		-- colors: 40, 40, 40, 40
			        8961 => x"00000000",		-- colors: 40, 40, 40, 40
			        8962 => x"00000000",		-- colors: 40, 40, 40, 40
			        8963 => x"00000000",		-- colors: 40, 40, 40, 40
			        8964 => x"00000000",		-- colors: 40, 40, 40, 40
			        8965 => x"00000000",		-- colors: 40, 40, 40, 40
			        8966 => x"00000000",		-- colors: 40, 40, 40, 40
			        8967 => x"00000000",		-- colors: 40, 40, 40, 40
			        8968 => x"00000000",		-- colors: 40, 40, 40, 40
			        8969 => x"00000000",		-- colors: 40, 40, 40, 40
			        8970 => x"00000000",		-- colors: 40, 40, 40, 40
			        8971 => x"00000000",		-- colors: 40, 40, 40, 40
			        8972 => x"00000000",		-- colors: 40, 40, 40, 40
			        8973 => x"00000000",		-- colors: 40, 40, 40, 40
			        8974 => x"00000000",		-- colors: 40, 40, 40, 40
			        8975 => x"00000000",		-- colors: 40, 40, 40, 40
			        8976 => x"00000000",		-- colors: 40, 40, 40, 40
			        8977 => x"00000000",		-- colors: 40, 40, 40, 40
			        8978 => x"00000000",		-- colors: 40, 40, 40, 40
			        8979 => x"00000000",		-- colors: 40, 40, 40, 40
			        8980 => x"00000000",		-- colors: 40, 40, 40, 40
			        8981 => x"00000000",		-- colors: 40, 40, 40, 40
			        8982 => x"00000000",		-- colors: 40, 40, 40, 40
			        8983 => x"00000000",		-- colors: 40, 40, 40, 40
			        8984 => x"00000000",		-- colors: 40, 40, 40, 40
			        8985 => x"00000000",		-- colors: 40, 40, 40, 40
			        8986 => x"00000000",		-- colors: 40, 40, 40, 40
			        8987 => x"00000000",		-- colors: 40, 40, 40, 40
			        8988 => x"00000000",		-- colors: 40, 40, 40, 40
			        8989 => x"00000000",		-- colors: 40, 40, 40, 40
			        8990 => x"00000000",		-- colors: 40, 40, 40, 40
			        8991 => x"00000000",		-- colors: 40, 40, 40, 40
			        8992 => x"00000000",		-- colors: 40, 40, 40, 40
			        8993 => x"00000000",		-- colors: 40, 40, 40, 40
			        8994 => x"00000000",		-- colors: 40, 40, 40, 40
			        8995 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8996 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8997 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8998 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        8999 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9000 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9001 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9002 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9003 => x"00000000",		-- colors: 40, 40, 40, 40
			        9004 => x"00000000",		-- colors: 40, 40, 40, 40
			        9005 => x"00000000",		-- colors: 40, 40, 40, 40
			        9006 => x"00000000",		-- colors: 40, 40, 40, 40
			        9007 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9008 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9009 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9010 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9011 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9012 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9013 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9014 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9015 => x"00000000",		-- colors: 40, 40, 40, 40
			        9016 => x"00000000",		-- colors: 40, 40, 40, 40
			        9017 => x"00000000",		-- colors: 40, 40, 40, 40
			        9018 => x"00000000",		-- colors: 40, 40, 40, 40
			        9019 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9020 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9021 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9022 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60

			                --  sprite 137
			        9023 => x"00000000",		-- colors: 40, 40, 40, 40
			        9024 => x"00000000",		-- colors: 40, 40, 40, 40
			        9025 => x"00000000",		-- colors: 40, 40, 40, 40
			        9026 => x"00000000",		-- colors: 40, 40, 40, 40
			        9027 => x"00000000",		-- colors: 40, 40, 40, 40
			        9028 => x"00000000",		-- colors: 40, 40, 40, 40
			        9029 => x"00000000",		-- colors: 40, 40, 40, 40
			        9030 => x"00000000",		-- colors: 40, 40, 40, 40
			        9031 => x"00000000",		-- colors: 40, 40, 40, 40
			        9032 => x"00000000",		-- colors: 40, 40, 40, 40
			        9033 => x"00000000",		-- colors: 40, 40, 40, 40
			        9034 => x"00000000",		-- colors: 40, 40, 40, 40
			        9035 => x"00000000",		-- colors: 40, 40, 40, 40
			        9036 => x"00000000",		-- colors: 40, 40, 40, 40
			        9037 => x"00000000",		-- colors: 40, 40, 40, 40
			        9038 => x"00000000",		-- colors: 40, 40, 40, 40
			        9039 => x"00000000",		-- colors: 40, 40, 40, 40
			        9040 => x"00000000",		-- colors: 40, 40, 40, 40
			        9041 => x"00000000",		-- colors: 40, 40, 40, 40
			        9042 => x"00000000",		-- colors: 40, 40, 40, 40
			        9043 => x"00000000",		-- colors: 40, 40, 40, 40
			        9044 => x"00000000",		-- colors: 40, 40, 40, 40
			        9045 => x"00000000",		-- colors: 40, 40, 40, 40
			        9046 => x"00000000",		-- colors: 40, 40, 40, 40
			        9047 => x"00000000",		-- colors: 40, 40, 40, 40
			        9048 => x"00000000",		-- colors: 40, 40, 40, 40
			        9049 => x"00000000",		-- colors: 40, 40, 40, 40
			        9050 => x"00000000",		-- colors: 40, 40, 40, 40
			        9051 => x"00000000",		-- colors: 40, 40, 40, 40
			        9052 => x"00000000",		-- colors: 40, 40, 40, 40
			        9053 => x"00000000",		-- colors: 40, 40, 40, 40
			        9054 => x"00000000",		-- colors: 40, 40, 40, 40
			        9055 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9056 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9057 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9058 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9059 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9060 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9061 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9062 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9063 => x"00000000",		-- colors: 40, 40, 40, 40
			        9064 => x"00000000",		-- colors: 40, 40, 40, 40
			        9065 => x"00000000",		-- colors: 40, 40, 40, 40
			        9066 => x"00000000",		-- colors: 40, 40, 40, 40
			        9067 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9068 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9069 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9070 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9071 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9072 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9073 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9074 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9075 => x"00000000",		-- colors: 40, 40, 40, 40
			        9076 => x"00000000",		-- colors: 40, 40, 40, 40
			        9077 => x"00000000",		-- colors: 40, 40, 40, 40
			        9078 => x"00000000",		-- colors: 40, 40, 40, 40
			        9079 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9080 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9081 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9082 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9083 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9084 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9085 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9086 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60

			                --  sprite 138
			        9087 => x"00000000",		-- colors: 40, 40, 40, 40
			        9088 => x"00000000",		-- colors: 40, 40, 40, 40
			        9089 => x"00000000",		-- colors: 40, 40, 40, 40
			        9090 => x"00000000",		-- colors: 40, 40, 40, 40
			        9091 => x"00000000",		-- colors: 40, 40, 40, 40
			        9092 => x"00000000",		-- colors: 40, 40, 40, 40
			        9093 => x"00000000",		-- colors: 40, 40, 40, 40
			        9094 => x"00000000",		-- colors: 40, 40, 40, 40
			        9095 => x"00000000",		-- colors: 40, 40, 40, 40
			        9096 => x"00000000",		-- colors: 40, 40, 40, 40
			        9097 => x"00000000",		-- colors: 40, 40, 40, 40
			        9098 => x"00000000",		-- colors: 40, 40, 40, 40
			        9099 => x"00000000",		-- colors: 40, 40, 40, 40
			        9100 => x"00000000",		-- colors: 40, 40, 40, 40
			        9101 => x"00000000",		-- colors: 40, 40, 40, 40
			        9102 => x"00000000",		-- colors: 40, 40, 40, 40
			        9103 => x"00000000",		-- colors: 40, 40, 40, 40
			        9104 => x"00000000",		-- colors: 40, 40, 40, 40
			        9105 => x"00000000",		-- colors: 40, 40, 40, 40
			        9106 => x"00000000",		-- colors: 40, 40, 40, 40
			        9107 => x"00000000",		-- colors: 40, 40, 40, 40
			        9108 => x"00000000",		-- colors: 40, 40, 40, 40
			        9109 => x"00000000",		-- colors: 40, 40, 40, 40
			        9110 => x"00000000",		-- colors: 40, 40, 40, 40
			        9111 => x"00000000",		-- colors: 40, 40, 40, 40
			        9112 => x"00000000",		-- colors: 40, 40, 40, 40
			        9113 => x"00000000",		-- colors: 40, 40, 40, 40
			        9114 => x"00000000",		-- colors: 40, 40, 40, 40
			        9115 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9116 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9117 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9118 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9119 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9120 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9121 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9122 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9123 => x"00000000",		-- colors: 40, 40, 40, 40
			        9124 => x"00000000",		-- colors: 40, 40, 40, 40
			        9125 => x"00000000",		-- colors: 40, 40, 40, 40
			        9126 => x"00000000",		-- colors: 40, 40, 40, 40
			        9127 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9128 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9129 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9130 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9131 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9132 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9133 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9134 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9135 => x"00000000",		-- colors: 40, 40, 40, 40
			        9136 => x"00000000",		-- colors: 40, 40, 40, 40
			        9137 => x"00000000",		-- colors: 40, 40, 40, 40
			        9138 => x"00000000",		-- colors: 40, 40, 40, 40
			        9139 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9140 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9141 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9142 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9143 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9144 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9145 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9146 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9147 => x"00000000",		-- colors: 40, 40, 40, 40
			        9148 => x"00000000",		-- colors: 40, 40, 40, 40
			        9149 => x"00000000",		-- colors: 40, 40, 40, 40
			        9150 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 139
			        9151 => x"00000000",		-- colors: 40, 40, 40, 40
			        9152 => x"00000000",		-- colors: 40, 40, 40, 40
			        9153 => x"00000000",		-- colors: 40, 40, 40, 40
			        9154 => x"00000000",		-- colors: 40, 40, 40, 40
			        9155 => x"00000000",		-- colors: 40, 40, 40, 40
			        9156 => x"00000000",		-- colors: 40, 40, 40, 40
			        9157 => x"00000000",		-- colors: 40, 40, 40, 40
			        9158 => x"00000000",		-- colors: 40, 40, 40, 40
			        9159 => x"00000000",		-- colors: 40, 40, 40, 40
			        9160 => x"00000000",		-- colors: 40, 40, 40, 40
			        9161 => x"00000000",		-- colors: 40, 40, 40, 40
			        9162 => x"00000000",		-- colors: 40, 40, 40, 40
			        9163 => x"00000000",		-- colors: 40, 40, 40, 40
			        9164 => x"00000000",		-- colors: 40, 40, 40, 40
			        9165 => x"00000000",		-- colors: 40, 40, 40, 40
			        9166 => x"00000000",		-- colors: 40, 40, 40, 40
			        9167 => x"00000000",		-- colors: 40, 40, 40, 40
			        9168 => x"00000000",		-- colors: 40, 40, 40, 40
			        9169 => x"00000000",		-- colors: 40, 40, 40, 40
			        9170 => x"00000000",		-- colors: 40, 40, 40, 40
			        9171 => x"00000000",		-- colors: 40, 40, 40, 40
			        9172 => x"00000000",		-- colors: 40, 40, 40, 40
			        9173 => x"00000000",		-- colors: 40, 40, 40, 40
			        9174 => x"00000000",		-- colors: 40, 40, 40, 40
			        9175 => x"00000000",		-- colors: 40, 40, 40, 40
			        9176 => x"00000000",		-- colors: 40, 40, 40, 40
			        9177 => x"00000000",		-- colors: 40, 40, 40, 40
			        9178 => x"00000000",		-- colors: 40, 40, 40, 40
			        9179 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9180 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9181 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9182 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9183 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9184 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9185 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9186 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9187 => x"00000000",		-- colors: 40, 40, 40, 40
			        9188 => x"00000000",		-- colors: 40, 40, 40, 40
			        9189 => x"00000000",		-- colors: 40, 40, 40, 40
			        9190 => x"00000000",		-- colors: 40, 40, 40, 40
			        9191 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9192 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9193 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9194 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9195 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9196 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9197 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9198 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9199 => x"00000000",		-- colors: 40, 40, 40, 40
			        9200 => x"00000000",		-- colors: 40, 40, 40, 40
			        9201 => x"00000000",		-- colors: 40, 40, 40, 40
			        9202 => x"00000000",		-- colors: 40, 40, 40, 40
			        9203 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9204 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9205 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9206 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9207 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9208 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9209 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9210 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9211 => x"00000000",		-- colors: 40, 40, 40, 40
			        9212 => x"00000000",		-- colors: 40, 40, 40, 40
			        9213 => x"00000000",		-- colors: 40, 40, 40, 40
			        9214 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 140
			        9215 => x"00000000",		-- colors: 40, 40, 40, 40
			        9216 => x"00000000",		-- colors: 40, 40, 40, 40
			        9217 => x"00000000",		-- colors: 40, 40, 40, 40
			        9218 => x"00000000",		-- colors: 40, 40, 40, 40
			        9219 => x"00000000",		-- colors: 40, 40, 40, 40
			        9220 => x"00000000",		-- colors: 40, 40, 40, 40
			        9221 => x"00000000",		-- colors: 40, 40, 40, 40
			        9222 => x"00000000",		-- colors: 40, 40, 40, 40
			        9223 => x"00000000",		-- colors: 40, 40, 40, 40
			        9224 => x"00000000",		-- colors: 40, 40, 40, 40
			        9225 => x"00000000",		-- colors: 40, 40, 40, 40
			        9226 => x"00000000",		-- colors: 40, 40, 40, 40
			        9227 => x"00000000",		-- colors: 40, 40, 40, 40
			        9228 => x"00000000",		-- colors: 40, 40, 40, 40
			        9229 => x"00000000",		-- colors: 40, 40, 40, 40
			        9230 => x"00000000",		-- colors: 40, 40, 40, 40
			        9231 => x"00000000",		-- colors: 40, 40, 40, 40
			        9232 => x"00000000",		-- colors: 40, 40, 40, 40
			        9233 => x"00000000",		-- colors: 40, 40, 40, 40
			        9234 => x"00000000",		-- colors: 40, 40, 40, 40
			        9235 => x"00000000",		-- colors: 40, 40, 40, 40
			        9236 => x"00000000",		-- colors: 40, 40, 40, 40
			        9237 => x"00000000",		-- colors: 40, 40, 40, 40
			        9238 => x"00000000",		-- colors: 40, 40, 40, 40
			        9239 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9240 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9241 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9242 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9243 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9244 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9245 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9246 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9247 => x"00000000",		-- colors: 40, 40, 40, 40
			        9248 => x"00000000",		-- colors: 40, 40, 40, 40
			        9249 => x"00000000",		-- colors: 40, 40, 40, 40
			        9250 => x"00000000",		-- colors: 40, 40, 40, 40
			        9251 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9252 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9253 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9254 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9255 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9256 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9257 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9258 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9259 => x"00000000",		-- colors: 40, 40, 40, 40
			        9260 => x"00000000",		-- colors: 40, 40, 40, 40
			        9261 => x"00000000",		-- colors: 40, 40, 40, 40
			        9262 => x"00000000",		-- colors: 40, 40, 40, 40
			        9263 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9264 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9265 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9266 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9267 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9268 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9269 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9270 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9271 => x"00000000",		-- colors: 40, 40, 40, 40
			        9272 => x"00000000",		-- colors: 40, 40, 40, 40
			        9273 => x"00000000",		-- colors: 40, 40, 40, 40
			        9274 => x"00000000",		-- colors: 40, 40, 40, 40
			        9275 => x"00000000",		-- colors: 40, 40, 40, 40
			        9276 => x"00000000",		-- colors: 40, 40, 40, 40
			        9277 => x"00000000",		-- colors: 40, 40, 40, 40
			        9278 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 141
			        9279 => x"00000000",		-- colors: 40, 40, 40, 40
			        9280 => x"00000000",		-- colors: 40, 40, 40, 40
			        9281 => x"00000000",		-- colors: 40, 40, 40, 40
			        9282 => x"00000000",		-- colors: 40, 40, 40, 40
			        9283 => x"00000000",		-- colors: 40, 40, 40, 40
			        9284 => x"00000000",		-- colors: 40, 40, 40, 40
			        9285 => x"00000000",		-- colors: 40, 40, 40, 40
			        9286 => x"00000000",		-- colors: 40, 40, 40, 40
			        9287 => x"32323232",		-- colors: 50, 50, 50, 50
			        9288 => x"32323232",		-- colors: 50, 50, 50, 50
			        9289 => x"32323232",		-- colors: 50, 50, 50, 50
			        9290 => x"32323232",		-- colors: 50, 50, 50, 50
			        9291 => x"00000000",		-- colors: 40, 40, 40, 40
			        9292 => x"00000000",		-- colors: 40, 40, 40, 40
			        9293 => x"00000000",		-- colors: 40, 40, 40, 40
			        9294 => x"00000000",		-- colors: 40, 40, 40, 40
			        9295 => x"00000000",		-- colors: 40, 40, 40, 40
			        9296 => x"00000000",		-- colors: 40, 40, 40, 40
			        9297 => x"00000000",		-- colors: 40, 40, 40, 40
			        9298 => x"00000000",		-- colors: 40, 40, 40, 40
			        9299 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9300 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9301 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9302 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9303 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9304 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9305 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9306 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9307 => x"00000000",		-- colors: 40, 40, 40, 40
			        9308 => x"00000000",		-- colors: 40, 40, 40, 40
			        9309 => x"00000000",		-- colors: 40, 40, 40, 40
			        9310 => x"00000000",		-- colors: 40, 40, 40, 40
			        9311 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9312 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9313 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9314 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9315 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9316 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9317 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9318 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9319 => x"00000000",		-- colors: 40, 40, 40, 40
			        9320 => x"00000000",		-- colors: 40, 40, 40, 40
			        9321 => x"00000000",		-- colors: 40, 40, 40, 40
			        9322 => x"00000000",		-- colors: 40, 40, 40, 40
			        9323 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9324 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9325 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9326 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9327 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9328 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9329 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9330 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9331 => x"00000000",		-- colors: 40, 40, 40, 40
			        9332 => x"00000000",		-- colors: 40, 40, 40, 40
			        9333 => x"00000000",		-- colors: 40, 40, 40, 40
			        9334 => x"00000000",		-- colors: 40, 40, 40, 40
			        9335 => x"00000000",		-- colors: 40, 40, 40, 40
			        9336 => x"00000000",		-- colors: 40, 40, 40, 40
			        9337 => x"00000000",		-- colors: 40, 40, 40, 40
			        9338 => x"00000000",		-- colors: 40, 40, 40, 40
			        9339 => x"00000000",		-- colors: 40, 40, 40, 40
			        9340 => x"00000000",		-- colors: 40, 40, 40, 40
			        9341 => x"00000000",		-- colors: 40, 40, 40, 40
			        9342 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 142
			        9343 => x"00000000",		-- colors: 40, 40, 40, 40
			        9344 => x"00000000",		-- colors: 40, 40, 40, 40
			        9345 => x"00000000",		-- colors: 40, 40, 40, 40
			        9346 => x"00000000",		-- colors: 40, 40, 40, 40
			        9347 => x"00000000",		-- colors: 40, 40, 40, 40
			        9348 => x"00000000",		-- colors: 40, 40, 40, 40
			        9349 => x"00000000",		-- colors: 40, 40, 40, 40
			        9350 => x"00000000",		-- colors: 40, 40, 40, 40
			        9351 => x"00000000",		-- colors: 40, 40, 40, 40
			        9352 => x"00000000",		-- colors: 40, 40, 40, 40
			        9353 => x"00000000",		-- colors: 40, 40, 40, 40
			        9354 => x"00000000",		-- colors: 40, 40, 40, 40
			        9355 => x"00000000",		-- colors: 40, 40, 40, 40
			        9356 => x"00000000",		-- colors: 40, 40, 40, 40
			        9357 => x"00000000",		-- colors: 40, 40, 40, 40
			        9358 => x"00000000",		-- colors: 40, 40, 40, 40
			        9359 => x"00000000",		-- colors: 40, 40, 40, 40
			        9360 => x"00000000",		-- colors: 40, 40, 40, 40
			        9361 => x"00000000",		-- colors: 40, 40, 40, 40
			        9362 => x"00000000",		-- colors: 40, 40, 40, 40
			        9363 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9364 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9365 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9366 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9367 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9368 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9369 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9370 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9371 => x"00000000",		-- colors: 40, 40, 40, 40
			        9372 => x"00000000",		-- colors: 40, 40, 40, 40
			        9373 => x"00000000",		-- colors: 40, 40, 40, 40
			        9374 => x"00000000",		-- colors: 40, 40, 40, 40
			        9375 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9376 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9377 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9378 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9379 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9380 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9381 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9382 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9383 => x"00000000",		-- colors: 40, 40, 40, 40
			        9384 => x"00000000",		-- colors: 40, 40, 40, 40
			        9385 => x"00000000",		-- colors: 40, 40, 40, 40
			        9386 => x"00000000",		-- colors: 40, 40, 40, 40
			        9387 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9388 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9389 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9390 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9391 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9392 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9393 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9394 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9395 => x"00000000",		-- colors: 40, 40, 40, 40
			        9396 => x"00000000",		-- colors: 40, 40, 40, 40
			        9397 => x"00000000",		-- colors: 40, 40, 40, 40
			        9398 => x"00000000",		-- colors: 40, 40, 40, 40
			        9399 => x"00000000",		-- colors: 40, 40, 40, 40
			        9400 => x"00000000",		-- colors: 40, 40, 40, 40
			        9401 => x"00000000",		-- colors: 40, 40, 40, 40
			        9402 => x"00000000",		-- colors: 40, 40, 40, 40
			        9403 => x"00000000",		-- colors: 40, 40, 40, 40
			        9404 => x"00000000",		-- colors: 40, 40, 40, 40
			        9405 => x"00000000",		-- colors: 40, 40, 40, 40
			        9406 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 143
			        9407 => x"00000000",		-- colors: 40, 40, 40, 40
			        9408 => x"00000000",		-- colors: 40, 40, 40, 40
			        9409 => x"00000000",		-- colors: 40, 40, 40, 40
			        9410 => x"00000000",		-- colors: 40, 40, 40, 40
			        9411 => x"00000000",		-- colors: 40, 40, 40, 40
			        9412 => x"00000000",		-- colors: 40, 40, 40, 40
			        9413 => x"00000000",		-- colors: 40, 40, 40, 40
			        9414 => x"00000000",		-- colors: 40, 40, 40, 40
			        9415 => x"00000000",		-- colors: 40, 40, 40, 40
			        9416 => x"00000000",		-- colors: 40, 40, 40, 40
			        9417 => x"00000000",		-- colors: 40, 40, 40, 40
			        9418 => x"00000000",		-- colors: 40, 40, 40, 40
			        9419 => x"00000000",		-- colors: 40, 40, 40, 40
			        9420 => x"00000000",		-- colors: 40, 40, 40, 40
			        9421 => x"00000000",		-- colors: 40, 40, 40, 40
			        9422 => x"00000000",		-- colors: 40, 40, 40, 40
			        9423 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9424 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9425 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9426 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9427 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9428 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9429 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9430 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9431 => x"00000000",		-- colors: 40, 40, 40, 40
			        9432 => x"00000000",		-- colors: 40, 40, 40, 40
			        9433 => x"00000000",		-- colors: 40, 40, 40, 40
			        9434 => x"00000000",		-- colors: 40, 40, 40, 40
			        9435 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9436 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9437 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9438 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9439 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9440 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9441 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9442 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9443 => x"00000000",		-- colors: 40, 40, 40, 40
			        9444 => x"00000000",		-- colors: 40, 40, 40, 40
			        9445 => x"00000000",		-- colors: 40, 40, 40, 40
			        9446 => x"00000000",		-- colors: 40, 40, 40, 40
			        9447 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9448 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9449 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9450 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9451 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9452 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9453 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9454 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9455 => x"00000000",		-- colors: 40, 40, 40, 40
			        9456 => x"00000000",		-- colors: 40, 40, 40, 40
			        9457 => x"00000000",		-- colors: 40, 40, 40, 40
			        9458 => x"00000000",		-- colors: 40, 40, 40, 40
			        9459 => x"00000000",		-- colors: 40, 40, 40, 40
			        9460 => x"00000000",		-- colors: 40, 40, 40, 40
			        9461 => x"00000000",		-- colors: 40, 40, 40, 40
			        9462 => x"00000000",		-- colors: 40, 40, 40, 40
			        9463 => x"00000000",		-- colors: 40, 40, 40, 40
			        9464 => x"00000000",		-- colors: 40, 40, 40, 40
			        9465 => x"00000000",		-- colors: 40, 40, 40, 40
			        9466 => x"00000000",		-- colors: 40, 40, 40, 40
			        9467 => x"00000000",		-- colors: 40, 40, 40, 40
			        9468 => x"00000000",		-- colors: 40, 40, 40, 40
			        9469 => x"00000000",		-- colors: 40, 40, 40, 40
			        9470 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 144
			        9471 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9472 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9473 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9474 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9475 => x"00000000",		-- colors: 40, 40, 40, 40
			        9476 => x"00000000",		-- colors: 40, 40, 40, 40
			        9477 => x"00000000",		-- colors: 40, 40, 40, 40
			        9478 => x"00000000",		-- colors: 40, 40, 40, 40
			        9479 => x"00000000",		-- colors: 40, 40, 40, 40
			        9480 => x"00000000",		-- colors: 40, 40, 40, 40
			        9481 => x"00000000",		-- colors: 40, 40, 40, 40
			        9482 => x"00000000",		-- colors: 40, 40, 40, 40
			        9483 => x"00000000",		-- colors: 40, 40, 40, 40
			        9484 => x"00000000",		-- colors: 40, 40, 40, 40
			        9485 => x"00000000",		-- colors: 40, 40, 40, 40
			        9486 => x"00000000",		-- colors: 40, 40, 40, 40
			        9487 => x"00000000",		-- colors: 40, 40, 40, 40
			        9488 => x"00000000",		-- colors: 40, 40, 40, 40
			        9489 => x"00000000",		-- colors: 40, 40, 40, 40
			        9490 => x"00000000",		-- colors: 40, 40, 40, 40
			        9491 => x"00000000",		-- colors: 40, 40, 40, 40
			        9492 => x"00000000",		-- colors: 40, 40, 40, 40
			        9493 => x"00000000",		-- colors: 40, 40, 40, 40
			        9494 => x"00000000",		-- colors: 40, 40, 40, 40
			        9495 => x"00000000",		-- colors: 40, 40, 40, 40
			        9496 => x"00000000",		-- colors: 40, 40, 40, 40
			        9497 => x"00000000",		-- colors: 40, 40, 40, 40
			        9498 => x"00000000",		-- colors: 40, 40, 40, 40
			        9499 => x"00000000",		-- colors: 40, 40, 40, 40
			        9500 => x"00000000",		-- colors: 40, 40, 40, 40
			        9501 => x"00000000",		-- colors: 40, 40, 40, 40
			        9502 => x"00000000",		-- colors: 40, 40, 40, 40
			        9503 => x"00000000",		-- colors: 40, 40, 40, 40
			        9504 => x"00000000",		-- colors: 40, 40, 40, 40
			        9505 => x"00000000",		-- colors: 40, 40, 40, 40
			        9506 => x"00000000",		-- colors: 40, 40, 40, 40
			        9507 => x"00000000",		-- colors: 40, 40, 40, 40
			        9508 => x"00000000",		-- colors: 40, 40, 40, 40
			        9509 => x"00000000",		-- colors: 40, 40, 40, 40
			        9510 => x"00000000",		-- colors: 40, 40, 40, 40
			        9511 => x"00000000",		-- colors: 40, 40, 40, 40
			        9512 => x"00000000",		-- colors: 40, 40, 40, 40
			        9513 => x"00000000",		-- colors: 40, 40, 40, 40
			        9514 => x"00000000",		-- colors: 40, 40, 40, 40
			        9515 => x"00000000",		-- colors: 40, 40, 40, 40
			        9516 => x"00000000",		-- colors: 40, 40, 40, 40
			        9517 => x"00000000",		-- colors: 40, 40, 40, 40
			        9518 => x"00000000",		-- colors: 40, 40, 40, 40
			        9519 => x"00000000",		-- colors: 40, 40, 40, 40
			        9520 => x"00000000",		-- colors: 40, 40, 40, 40
			        9521 => x"00000000",		-- colors: 40, 40, 40, 40
			        9522 => x"00000000",		-- colors: 40, 40, 40, 40
			        9523 => x"00000000",		-- colors: 40, 40, 40, 40
			        9524 => x"00000000",		-- colors: 40, 40, 40, 40
			        9525 => x"00000000",		-- colors: 40, 40, 40, 40
			        9526 => x"00000000",		-- colors: 40, 40, 40, 40
			        9527 => x"00000000",		-- colors: 40, 40, 40, 40
			        9528 => x"00000000",		-- colors: 40, 40, 40, 40
			        9529 => x"00000000",		-- colors: 40, 40, 40, 40
			        9530 => x"00000000",		-- colors: 40, 40, 40, 40
			        9531 => x"00000000",		-- colors: 40, 40, 40, 40
			        9532 => x"00000000",		-- colors: 40, 40, 40, 40
			        9533 => x"00000000",		-- colors: 40, 40, 40, 40
			        9534 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 145
			        9535 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9536 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9537 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9538 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9539 => x"00000000",		-- colors: 40, 40, 40, 40
			        9540 => x"00000000",		-- colors: 40, 40, 40, 40
			        9541 => x"00000000",		-- colors: 40, 40, 40, 40
			        9542 => x"00000000",		-- colors: 40, 40, 40, 40
			        9543 => x"00000000",		-- colors: 40, 40, 40, 40
			        9544 => x"00000000",		-- colors: 40, 40, 40, 40
			        9545 => x"00000000",		-- colors: 40, 40, 40, 40
			        9546 => x"00000000",		-- colors: 40, 40, 40, 40
			        9547 => x"00000000",		-- colors: 40, 40, 40, 40
			        9548 => x"00000000",		-- colors: 40, 40, 40, 40
			        9549 => x"00000000",		-- colors: 40, 40, 40, 40
			        9550 => x"00000000",		-- colors: 40, 40, 40, 40
			        9551 => x"00000000",		-- colors: 40, 40, 40, 40
			        9552 => x"00000000",		-- colors: 40, 40, 40, 40
			        9553 => x"00000000",		-- colors: 40, 40, 40, 40
			        9554 => x"00000000",		-- colors: 40, 40, 40, 40
			        9555 => x"00000000",		-- colors: 40, 40, 40, 40
			        9556 => x"00000000",		-- colors: 40, 40, 40, 40
			        9557 => x"00000000",		-- colors: 40, 40, 40, 40
			        9558 => x"00000000",		-- colors: 40, 40, 40, 40
			        9559 => x"00000000",		-- colors: 40, 40, 40, 40
			        9560 => x"00000000",		-- colors: 40, 40, 40, 40
			        9561 => x"00000000",		-- colors: 40, 40, 40, 40
			        9562 => x"00000000",		-- colors: 40, 40, 40, 40
			        9563 => x"00000000",		-- colors: 40, 40, 40, 40
			        9564 => x"00000000",		-- colors: 40, 40, 40, 40
			        9565 => x"00000000",		-- colors: 40, 40, 40, 40
			        9566 => x"00000000",		-- colors: 40, 40, 40, 40
			        9567 => x"00000000",		-- colors: 40, 40, 40, 40
			        9568 => x"00000000",		-- colors: 40, 40, 40, 40
			        9569 => x"00000000",		-- colors: 40, 40, 40, 40
			        9570 => x"00000000",		-- colors: 40, 40, 40, 40
			        9571 => x"00000000",		-- colors: 40, 40, 40, 40
			        9572 => x"00000000",		-- colors: 40, 40, 40, 40
			        9573 => x"00000000",		-- colors: 40, 40, 40, 40
			        9574 => x"00000000",		-- colors: 40, 40, 40, 40
			        9575 => x"00000000",		-- colors: 40, 40, 40, 40
			        9576 => x"00000000",		-- colors: 40, 40, 40, 40
			        9577 => x"00000000",		-- colors: 40, 40, 40, 40
			        9578 => x"00000000",		-- colors: 40, 40, 40, 40
			        9579 => x"00000000",		-- colors: 40, 40, 40, 40
			        9580 => x"00000000",		-- colors: 40, 40, 40, 40
			        9581 => x"00000000",		-- colors: 40, 40, 40, 40
			        9582 => x"00000000",		-- colors: 40, 40, 40, 40
			        9583 => x"00000000",		-- colors: 40, 40, 40, 40
			        9584 => x"00000000",		-- colors: 40, 40, 40, 40
			        9585 => x"00000000",		-- colors: 40, 40, 40, 40
			        9586 => x"00000000",		-- colors: 40, 40, 40, 40
			        9587 => x"00000000",		-- colors: 40, 40, 40, 40
			        9588 => x"00000000",		-- colors: 40, 40, 40, 40
			        9589 => x"00000000",		-- colors: 40, 40, 40, 40
			        9590 => x"00000000",		-- colors: 40, 40, 40, 40
			        9591 => x"00000000",		-- colors: 40, 40, 40, 40
			        9592 => x"00000000",		-- colors: 40, 40, 40, 40
			        9593 => x"00000000",		-- colors: 40, 40, 40, 40
			        9594 => x"00000000",		-- colors: 40, 40, 40, 40
			        9595 => x"00000000",		-- colors: 40, 40, 40, 40
			        9596 => x"00000000",		-- colors: 40, 40, 40, 40
			        9597 => x"00000000",		-- colors: 40, 40, 40, 40
			        9598 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 146
			        9599 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9600 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9601 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9602 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9603 => x"00000000",		-- colors: 40, 40, 40, 40
			        9604 => x"00000000",		-- colors: 40, 40, 40, 40
			        9605 => x"00000000",		-- colors: 40, 40, 40, 40
			        9606 => x"00000000",		-- colors: 40, 40, 40, 40
			        9607 => x"00000000",		-- colors: 40, 40, 40, 40
			        9608 => x"00000000",		-- colors: 40, 40, 40, 40
			        9609 => x"00000000",		-- colors: 40, 40, 40, 40
			        9610 => x"00000000",		-- colors: 40, 40, 40, 40
			        9611 => x"00000000",		-- colors: 40, 40, 40, 40
			        9612 => x"00000000",		-- colors: 40, 40, 40, 40
			        9613 => x"00000000",		-- colors: 40, 40, 40, 40
			        9614 => x"00000000",		-- colors: 40, 40, 40, 40
			        9615 => x"00000000",		-- colors: 40, 40, 40, 40
			        9616 => x"00000000",		-- colors: 40, 40, 40, 40
			        9617 => x"00000000",		-- colors: 40, 40, 40, 40
			        9618 => x"00000000",		-- colors: 40, 40, 40, 40
			        9619 => x"00000000",		-- colors: 40, 40, 40, 40
			        9620 => x"00000000",		-- colors: 40, 40, 40, 40
			        9621 => x"00000000",		-- colors: 40, 40, 40, 40
			        9622 => x"00000000",		-- colors: 40, 40, 40, 40
			        9623 => x"00000000",		-- colors: 40, 40, 40, 40
			        9624 => x"00000000",		-- colors: 40, 40, 40, 40
			        9625 => x"00000000",		-- colors: 40, 40, 40, 40
			        9626 => x"00000000",		-- colors: 40, 40, 40, 40
			        9627 => x"00000000",		-- colors: 40, 40, 40, 40
			        9628 => x"00000000",		-- colors: 40, 40, 40, 40
			        9629 => x"00000000",		-- colors: 40, 40, 40, 40
			        9630 => x"00000000",		-- colors: 40, 40, 40, 40
			        9631 => x"00000000",		-- colors: 40, 40, 40, 40
			        9632 => x"00000000",		-- colors: 40, 40, 40, 40
			        9633 => x"00000000",		-- colors: 40, 40, 40, 40
			        9634 => x"00000000",		-- colors: 40, 40, 40, 40
			        9635 => x"00000000",		-- colors: 40, 40, 40, 40
			        9636 => x"00000000",		-- colors: 40, 40, 40, 40
			        9637 => x"00000000",		-- colors: 40, 40, 40, 40
			        9638 => x"00000000",		-- colors: 40, 40, 40, 40
			        9639 => x"00000000",		-- colors: 40, 40, 40, 40
			        9640 => x"00000000",		-- colors: 40, 40, 40, 40
			        9641 => x"00000000",		-- colors: 40, 40, 40, 40
			        9642 => x"00000000",		-- colors: 40, 40, 40, 40
			        9643 => x"00000000",		-- colors: 40, 40, 40, 40
			        9644 => x"00000000",		-- colors: 40, 40, 40, 40
			        9645 => x"00000000",		-- colors: 40, 40, 40, 40
			        9646 => x"00000000",		-- colors: 40, 40, 40, 40
			        9647 => x"00000000",		-- colors: 40, 40, 40, 40
			        9648 => x"00000000",		-- colors: 40, 40, 40, 40
			        9649 => x"00000000",		-- colors: 40, 40, 40, 40
			        9650 => x"00000000",		-- colors: 40, 40, 40, 40
			        9651 => x"00000000",		-- colors: 40, 40, 40, 40
			        9652 => x"00000000",		-- colors: 40, 40, 40, 40
			        9653 => x"00000000",		-- colors: 40, 40, 40, 40
			        9654 => x"00000000",		-- colors: 40, 40, 40, 40
			        9655 => x"00000000",		-- colors: 40, 40, 40, 40
			        9656 => x"00000000",		-- colors: 40, 40, 40, 40
			        9657 => x"00000000",		-- colors: 40, 40, 40, 40
			        9658 => x"00000000",		-- colors: 40, 40, 40, 40
			        9659 => x"00000000",		-- colors: 40, 40, 40, 40
			        9660 => x"00000000",		-- colors: 40, 40, 40, 40
			        9661 => x"00000000",		-- colors: 40, 40, 40, 40
			        9662 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 147
			        9663 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9664 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9665 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9666 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9667 => x"00000000",		-- colors: 40, 40, 40, 40
			        9668 => x"00000000",		-- colors: 40, 40, 40, 40
			        9669 => x"00000000",		-- colors: 40, 40, 40, 40
			        9670 => x"00000000",		-- colors: 40, 40, 40, 40
			        9671 => x"00000000",		-- colors: 40, 40, 40, 40
			        9672 => x"00000000",		-- colors: 40, 40, 40, 40
			        9673 => x"00000000",		-- colors: 40, 40, 40, 40
			        9674 => x"00000000",		-- colors: 40, 40, 40, 40
			        9675 => x"00000000",		-- colors: 40, 40, 40, 40
			        9676 => x"00000000",		-- colors: 40, 40, 40, 40
			        9677 => x"00000000",		-- colors: 40, 40, 40, 40
			        9678 => x"00000000",		-- colors: 40, 40, 40, 40
			        9679 => x"00000000",		-- colors: 40, 40, 40, 40
			        9680 => x"00000000",		-- colors: 40, 40, 40, 40
			        9681 => x"00000000",		-- colors: 40, 40, 40, 40
			        9682 => x"00000000",		-- colors: 40, 40, 40, 40
			        9683 => x"00000000",		-- colors: 40, 40, 40, 40
			        9684 => x"00000000",		-- colors: 40, 40, 40, 40
			        9685 => x"00000000",		-- colors: 40, 40, 40, 40
			        9686 => x"00000000",		-- colors: 40, 40, 40, 40
			        9687 => x"00000000",		-- colors: 40, 40, 40, 40
			        9688 => x"00000000",		-- colors: 40, 40, 40, 40
			        9689 => x"00000000",		-- colors: 40, 40, 40, 40
			        9690 => x"00000000",		-- colors: 40, 40, 40, 40
			        9691 => x"00000000",		-- colors: 40, 40, 40, 40
			        9692 => x"00000000",		-- colors: 40, 40, 40, 40
			        9693 => x"00000000",		-- colors: 40, 40, 40, 40
			        9694 => x"00000000",		-- colors: 40, 40, 40, 40
			        9695 => x"00000000",		-- colors: 40, 40, 40, 40
			        9696 => x"00000000",		-- colors: 40, 40, 40, 40
			        9697 => x"00000000",		-- colors: 40, 40, 40, 40
			        9698 => x"00000000",		-- colors: 40, 40, 40, 40
			        9699 => x"00000000",		-- colors: 40, 40, 40, 40
			        9700 => x"00000000",		-- colors: 40, 40, 40, 40
			        9701 => x"00000000",		-- colors: 40, 40, 40, 40
			        9702 => x"00000000",		-- colors: 40, 40, 40, 40
			        9703 => x"00000000",		-- colors: 40, 40, 40, 40
			        9704 => x"00000000",		-- colors: 40, 40, 40, 40
			        9705 => x"00000000",		-- colors: 40, 40, 40, 40
			        9706 => x"00000000",		-- colors: 40, 40, 40, 40
			        9707 => x"00000000",		-- colors: 40, 40, 40, 40
			        9708 => x"00000000",		-- colors: 40, 40, 40, 40
			        9709 => x"00000000",		-- colors: 40, 40, 40, 40
			        9710 => x"00000000",		-- colors: 40, 40, 40, 40
			        9711 => x"00000000",		-- colors: 40, 40, 40, 40
			        9712 => x"00000000",		-- colors: 40, 40, 40, 40
			        9713 => x"00000000",		-- colors: 40, 40, 40, 40
			        9714 => x"00000000",		-- colors: 40, 40, 40, 40
			        9715 => x"00000000",		-- colors: 40, 40, 40, 40
			        9716 => x"00000000",		-- colors: 40, 40, 40, 40
			        9717 => x"00000000",		-- colors: 40, 40, 40, 40
			        9718 => x"00000000",		-- colors: 40, 40, 40, 40
			        9719 => x"00000000",		-- colors: 40, 40, 40, 40
			        9720 => x"00000000",		-- colors: 40, 40, 40, 40
			        9721 => x"00000000",		-- colors: 40, 40, 40, 40
			        9722 => x"00000000",		-- colors: 40, 40, 40, 40
			        9723 => x"00000000",		-- colors: 40, 40, 40, 40
			        9724 => x"00000000",		-- colors: 40, 40, 40, 40
			        9725 => x"00000000",		-- colors: 40, 40, 40, 40
			        9726 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 148
			        9727 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9728 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9729 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9730 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9731 => x"00000000",		-- colors: 40, 40, 40, 40
			        9732 => x"00000000",		-- colors: 40, 40, 40, 40
			        9733 => x"00000000",		-- colors: 40, 40, 40, 40
			        9734 => x"00000000",		-- colors: 40, 40, 40, 40
			        9735 => x"00000000",		-- colors: 40, 40, 40, 40
			        9736 => x"00000000",		-- colors: 40, 40, 40, 40
			        9737 => x"00000000",		-- colors: 40, 40, 40, 40
			        9738 => x"00000000",		-- colors: 40, 40, 40, 40
			        9739 => x"00000000",		-- colors: 40, 40, 40, 40
			        9740 => x"00000000",		-- colors: 40, 40, 40, 40
			        9741 => x"00000000",		-- colors: 40, 40, 40, 40
			        9742 => x"00000000",		-- colors: 40, 40, 40, 40
			        9743 => x"00000000",		-- colors: 40, 40, 40, 40
			        9744 => x"00000000",		-- colors: 40, 40, 40, 40
			        9745 => x"00000000",		-- colors: 40, 40, 40, 40
			        9746 => x"00000000",		-- colors: 40, 40, 40, 40
			        9747 => x"00000000",		-- colors: 40, 40, 40, 40
			        9748 => x"00000000",		-- colors: 40, 40, 40, 40
			        9749 => x"00000000",		-- colors: 40, 40, 40, 40
			        9750 => x"00000000",		-- colors: 40, 40, 40, 40
			        9751 => x"00000000",		-- colors: 40, 40, 40, 40
			        9752 => x"00000000",		-- colors: 40, 40, 40, 40
			        9753 => x"00000000",		-- colors: 40, 40, 40, 40
			        9754 => x"00000000",		-- colors: 40, 40, 40, 40
			        9755 => x"00000000",		-- colors: 40, 40, 40, 40
			        9756 => x"00000000",		-- colors: 40, 40, 40, 40
			        9757 => x"00000000",		-- colors: 40, 40, 40, 40
			        9758 => x"00000000",		-- colors: 40, 40, 40, 40
			        9759 => x"00000000",		-- colors: 40, 40, 40, 40
			        9760 => x"00000000",		-- colors: 40, 40, 40, 40
			        9761 => x"00000000",		-- colors: 40, 40, 40, 40
			        9762 => x"00000000",		-- colors: 40, 40, 40, 40
			        9763 => x"00000000",		-- colors: 40, 40, 40, 40
			        9764 => x"00000000",		-- colors: 40, 40, 40, 40
			        9765 => x"00000000",		-- colors: 40, 40, 40, 40
			        9766 => x"00000000",		-- colors: 40, 40, 40, 40
			        9767 => x"00000000",		-- colors: 40, 40, 40, 40
			        9768 => x"00000000",		-- colors: 40, 40, 40, 40
			        9769 => x"00000000",		-- colors: 40, 40, 40, 40
			        9770 => x"00000000",		-- colors: 40, 40, 40, 40
			        9771 => x"00000000",		-- colors: 40, 40, 40, 40
			        9772 => x"00000000",		-- colors: 40, 40, 40, 40
			        9773 => x"00000000",		-- colors: 40, 40, 40, 40
			        9774 => x"00000000",		-- colors: 40, 40, 40, 40
			        9775 => x"00000000",		-- colors: 40, 40, 40, 40
			        9776 => x"00000000",		-- colors: 40, 40, 40, 40
			        9777 => x"00000000",		-- colors: 40, 40, 40, 40
			        9778 => x"00000000",		-- colors: 40, 40, 40, 40
			        9779 => x"00000000",		-- colors: 40, 40, 40, 40
			        9780 => x"00000000",		-- colors: 40, 40, 40, 40
			        9781 => x"00000000",		-- colors: 40, 40, 40, 40
			        9782 => x"00000000",		-- colors: 40, 40, 40, 40
			        9783 => x"00000000",		-- colors: 40, 40, 40, 40
			        9784 => x"00000000",		-- colors: 40, 40, 40, 40
			        9785 => x"00000000",		-- colors: 40, 40, 40, 40
			        9786 => x"00000000",		-- colors: 40, 40, 40, 40
			        9787 => x"00000000",		-- colors: 40, 40, 40, 40
			        9788 => x"00000000",		-- colors: 40, 40, 40, 40
			        9789 => x"00000000",		-- colors: 40, 40, 40, 40
			        9790 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 149
			        9791 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9792 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9793 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9794 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9795 => x"00000000",		-- colors: 40, 40, 40, 40
			        9796 => x"00000000",		-- colors: 40, 40, 40, 40
			        9797 => x"00000000",		-- colors: 40, 40, 40, 40
			        9798 => x"00000000",		-- colors: 40, 40, 40, 40
			        9799 => x"00000000",		-- colors: 40, 40, 40, 40
			        9800 => x"00000000",		-- colors: 40, 40, 40, 40
			        9801 => x"00000000",		-- colors: 40, 40, 40, 40
			        9802 => x"00000000",		-- colors: 40, 40, 40, 40
			        9803 => x"00000000",		-- colors: 40, 40, 40, 40
			        9804 => x"00000000",		-- colors: 40, 40, 40, 40
			        9805 => x"00000000",		-- colors: 40, 40, 40, 40
			        9806 => x"00000000",		-- colors: 40, 40, 40, 40
			        9807 => x"00000000",		-- colors: 40, 40, 40, 40
			        9808 => x"00000000",		-- colors: 40, 40, 40, 40
			        9809 => x"00000000",		-- colors: 40, 40, 40, 40
			        9810 => x"00000000",		-- colors: 40, 40, 40, 40
			        9811 => x"00000000",		-- colors: 40, 40, 40, 40
			        9812 => x"00000000",		-- colors: 40, 40, 40, 40
			        9813 => x"00000000",		-- colors: 40, 40, 40, 40
			        9814 => x"00000000",		-- colors: 40, 40, 40, 40
			        9815 => x"00000000",		-- colors: 40, 40, 40, 40
			        9816 => x"00000000",		-- colors: 40, 40, 40, 40
			        9817 => x"00000000",		-- colors: 40, 40, 40, 40
			        9818 => x"00000000",		-- colors: 40, 40, 40, 40
			        9819 => x"00000000",		-- colors: 40, 40, 40, 40
			        9820 => x"00000000",		-- colors: 40, 40, 40, 40
			        9821 => x"00000000",		-- colors: 40, 40, 40, 40
			        9822 => x"00000000",		-- colors: 40, 40, 40, 40
			        9823 => x"00000000",		-- colors: 40, 40, 40, 40
			        9824 => x"00000000",		-- colors: 40, 40, 40, 40
			        9825 => x"00000000",		-- colors: 40, 40, 40, 40
			        9826 => x"00000000",		-- colors: 40, 40, 40, 40
			        9827 => x"00000000",		-- colors: 40, 40, 40, 40
			        9828 => x"00000000",		-- colors: 40, 40, 40, 40
			        9829 => x"00000000",		-- colors: 40, 40, 40, 40
			        9830 => x"00000000",		-- colors: 40, 40, 40, 40
			        9831 => x"00000000",		-- colors: 40, 40, 40, 40
			        9832 => x"00000000",		-- colors: 40, 40, 40, 40
			        9833 => x"00000000",		-- colors: 40, 40, 40, 40
			        9834 => x"00000000",		-- colors: 40, 40, 40, 40
			        9835 => x"00000000",		-- colors: 40, 40, 40, 40
			        9836 => x"00000000",		-- colors: 40, 40, 40, 40
			        9837 => x"00000000",		-- colors: 40, 40, 40, 40
			        9838 => x"00000000",		-- colors: 40, 40, 40, 40
			        9839 => x"00000000",		-- colors: 40, 40, 40, 40
			        9840 => x"00000000",		-- colors: 40, 40, 40, 40
			        9841 => x"00000000",		-- colors: 40, 40, 40, 40
			        9842 => x"00000000",		-- colors: 40, 40, 40, 40
			        9843 => x"00000000",		-- colors: 40, 40, 40, 40
			        9844 => x"00000000",		-- colors: 40, 40, 40, 40
			        9845 => x"00000000",		-- colors: 40, 40, 40, 40
			        9846 => x"00000000",		-- colors: 40, 40, 40, 40
			        9847 => x"00000000",		-- colors: 40, 40, 40, 40
			        9848 => x"00000000",		-- colors: 40, 40, 40, 40
			        9849 => x"00000000",		-- colors: 40, 40, 40, 40
			        9850 => x"00000000",		-- colors: 40, 40, 40, 40
			        9851 => x"00000000",		-- colors: 40, 40, 40, 40
			        9852 => x"00000000",		-- colors: 40, 40, 40, 40
			        9853 => x"00000000",		-- colors: 40, 40, 40, 40
			        9854 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 150
			        9855 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9856 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9857 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9858 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9859 => x"00000000",		-- colors: 40, 40, 40, 40
			        9860 => x"00000000",		-- colors: 40, 40, 40, 40
			        9861 => x"00000000",		-- colors: 40, 40, 40, 40
			        9862 => x"00000000",		-- colors: 40, 40, 40, 40
			        9863 => x"00000000",		-- colors: 40, 40, 40, 40
			        9864 => x"00000000",		-- colors: 40, 40, 40, 40
			        9865 => x"00000000",		-- colors: 40, 40, 40, 40
			        9866 => x"00000000",		-- colors: 40, 40, 40, 40
			        9867 => x"00000000",		-- colors: 40, 40, 40, 40
			        9868 => x"00000000",		-- colors: 40, 40, 40, 40
			        9869 => x"00000000",		-- colors: 40, 40, 40, 40
			        9870 => x"00000000",		-- colors: 40, 40, 40, 40
			        9871 => x"00000000",		-- colors: 40, 40, 40, 40
			        9872 => x"00000000",		-- colors: 40, 40, 40, 40
			        9873 => x"00000000",		-- colors: 40, 40, 40, 40
			        9874 => x"00000000",		-- colors: 40, 40, 40, 40
			        9875 => x"00000000",		-- colors: 40, 40, 40, 40
			        9876 => x"00000000",		-- colors: 40, 40, 40, 40
			        9877 => x"00000000",		-- colors: 40, 40, 40, 40
			        9878 => x"00000000",		-- colors: 40, 40, 40, 40
			        9879 => x"00000000",		-- colors: 40, 40, 40, 40
			        9880 => x"00000000",		-- colors: 40, 40, 40, 40
			        9881 => x"00000000",		-- colors: 40, 40, 40, 40
			        9882 => x"00000000",		-- colors: 40, 40, 40, 40
			        9883 => x"00000000",		-- colors: 40, 40, 40, 40
			        9884 => x"00000000",		-- colors: 40, 40, 40, 40
			        9885 => x"00000000",		-- colors: 40, 40, 40, 40
			        9886 => x"00000000",		-- colors: 40, 40, 40, 40
			        9887 => x"00000000",		-- colors: 40, 40, 40, 40
			        9888 => x"00000000",		-- colors: 40, 40, 40, 40
			        9889 => x"00000000",		-- colors: 40, 40, 40, 40
			        9890 => x"00000000",		-- colors: 40, 40, 40, 40
			        9891 => x"00000000",		-- colors: 40, 40, 40, 40
			        9892 => x"00000000",		-- colors: 40, 40, 40, 40
			        9893 => x"00000000",		-- colors: 40, 40, 40, 40
			        9894 => x"00000000",		-- colors: 40, 40, 40, 40
			        9895 => x"00000000",		-- colors: 40, 40, 40, 40
			        9896 => x"00000000",		-- colors: 40, 40, 40, 40
			        9897 => x"00000000",		-- colors: 40, 40, 40, 40
			        9898 => x"00000000",		-- colors: 40, 40, 40, 40
			        9899 => x"00000000",		-- colors: 40, 40, 40, 40
			        9900 => x"00000000",		-- colors: 40, 40, 40, 40
			        9901 => x"00000000",		-- colors: 40, 40, 40, 40
			        9902 => x"00000000",		-- colors: 40, 40, 40, 40
			        9903 => x"00000000",		-- colors: 40, 40, 40, 40
			        9904 => x"00000000",		-- colors: 40, 40, 40, 40
			        9905 => x"00000000",		-- colors: 40, 40, 40, 40
			        9906 => x"00000000",		-- colors: 40, 40, 40, 40
			        9907 => x"00000000",		-- colors: 40, 40, 40, 40
			        9908 => x"00000000",		-- colors: 40, 40, 40, 40
			        9909 => x"00000000",		-- colors: 40, 40, 40, 40
			        9910 => x"00000000",		-- colors: 40, 40, 40, 40
			        9911 => x"00000000",		-- colors: 40, 40, 40, 40
			        9912 => x"00000000",		-- colors: 40, 40, 40, 40
			        9913 => x"00000000",		-- colors: 40, 40, 40, 40
			        9914 => x"00000000",		-- colors: 40, 40, 40, 40
			        9915 => x"00000000",		-- colors: 40, 40, 40, 40
			        9916 => x"00000000",		-- colors: 40, 40, 40, 40
			        9917 => x"00000000",		-- colors: 40, 40, 40, 40
			        9918 => x"00000000",		-- colors: 40, 40, 40, 40

			                --  sprite 151
			        9919 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9920 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9921 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9922 => x"3C3C3C3C",		-- colors: 60, 60, 60, 60
			        9923 => x"00000000",		-- colors: 40, 40, 40, 40
			        9924 => x"00000000",		-- colors: 40, 40, 40, 40
			        9925 => x"00000000",		-- colors: 40, 40, 40, 40
			        9926 => x"00000000",		-- colors: 40, 40, 40, 40
			        9927 => x"00000000",		-- colors: 40, 40, 40, 40
			        9928 => x"00000000",		-- colors: 40, 40, 40, 40
			        9929 => x"00000000",		-- colors: 40, 40, 40, 40
			        9930 => x"00000000",		-- colors: 40, 40, 40, 40
			        9931 => x"00000000",		-- colors: 40, 40, 40, 40
			        9932 => x"00000000",		-- colors: 40, 40, 40, 40
			        9933 => x"00000000",		-- colors: 40, 40, 40, 40
			        9934 => x"00000000",		-- colors: 40, 40, 40, 40
			        9935 => x"00000000",		-- colors: 40, 40, 40, 40
			        9936 => x"00000000",		-- colors: 40, 40, 40, 40
			        9937 => x"00000000",		-- colors: 40, 40, 40, 40
			        9938 => x"00000000",		-- colors: 40, 40, 40, 40
			        9939 => x"00000000",		-- colors: 40, 40, 40, 40
			        9940 => x"00000000",		-- colors: 40, 40, 40, 40
			        9941 => x"00000000",		-- colors: 40, 40, 40, 40
			        9942 => x"00000000",		-- colors: 40, 40, 40, 40
			        9943 => x"00000000",		-- colors: 40, 40, 40, 40
			        9944 => x"00000000",		-- colors: 40, 40, 40, 40
			        9945 => x"00000000",		-- colors: 40, 40, 40, 40
			        9946 => x"00000000",		-- colors: 40, 40, 40, 40
			        9947 => x"00000000",		-- colors: 40, 40, 40, 40
			        9948 => x"00000000",		-- colors: 40, 40, 40, 40
			        9949 => x"00000000",		-- colors: 40, 40, 40, 40
			        9950 => x"00000000",		-- colors: 40, 40, 40, 40
			        9951 => x"00000000",		-- colors: 40, 40, 40, 40
			        9952 => x"00000000",		-- colors: 40, 40, 40, 40
			        9953 => x"00000000",		-- colors: 40, 40, 40, 40
			        9954 => x"00000000",		-- colors: 40, 40, 40, 40
			        9955 => x"00000000",		-- colors: 40, 40, 40, 40
			        9956 => x"00000000",		-- colors: 40, 40, 40, 40
			        9957 => x"00000000",		-- colors: 40, 40, 40, 40
			        9958 => x"00000000",		-- colors: 40, 40, 40, 40
			        9959 => x"00000000",		-- colors: 40, 40, 40, 40
			        9960 => x"00000000",		-- colors: 40, 40, 40, 40
			        9961 => x"00000000",		-- colors: 40, 40, 40, 40
			        9962 => x"00000000",		-- colors: 40, 40, 40, 40
			        9963 => x"00000000",		-- colors: 40, 40, 40, 40
			        9964 => x"00000000",		-- colors: 40, 40, 40, 40
			        9965 => x"00000000",		-- colors: 40, 40, 40, 40
			        9966 => x"00000000",		-- colors: 40, 40, 40, 40
			        9967 => x"00000000",		-- colors: 40, 40, 40, 40
			        9968 => x"00000000",		-- colors: 40, 40, 40, 40
			        9969 => x"00000000",		-- colors: 40, 40, 40, 40
			        9970 => x"00000000",		-- colors: 40, 40, 40, 40
			        9971 => x"00000000",		-- colors: 40, 40, 40, 40
			        9972 => x"00000000",		-- colors: 40, 40, 40, 40
			        9973 => x"00000000",		-- colors: 40, 40, 40, 40
			        9974 => x"00000000",		-- colors: 40, 40, 40, 40
			        9975 => x"00000000",		-- colors: 40, 40, 40, 40
			        9976 => x"00000000",		-- colors: 40, 40, 40, 40
			        9977 => x"00000000",		-- colors: 40, 40, 40, 40
			        9978 => x"00000000",		-- colors: 40, 40, 40, 40
			        9979 => x"00000000",		-- colors: 40, 40, 40, 40
			        9980 => x"00000000",		-- colors: 40, 40, 40, 40
			        9981 => x"00000000",		-- colors: 40, 40, 40, 40
			        9982 => x"00000000",		-- colors: 40, 40, 40, 40

				--		****  MAP  ****
				9983 => x"00000016", --padding
				9984 => x"00000016", --padding
				9985 => x"00000016", --padding
				9986 => x"00000016", --padding
				9987 => x"00000016", --padding
				9988 => x"00000016", --padding
				9989 => x"00000016", --padding
				9990 => x"00000016", --padding
				9991 => x"00000016", --padding
				9992 => x"00000016", --padding
				9993 => x"00000016", --padding
				9994 => x"00000016", --padding
				9995 => x"00000016", --padding
				9996 => x"00000016", --padding
				9997 => x"00000016", --padding
				9998 => x"00000016", --padding
				9999 => x"00000016", --padding
				10000 => x"00000016", --padding
				10001 => x"00000016", --padding
				10002 => x"00000016", --padding
				10003 => x"00000016", --padding
				10004 => x"00000016", --padding
				10005 => x"00000016", --padding
				10006 => x"00000016", --padding
				10007 => x"00000016", --padding
				10008 => x"00000016", --padding
				10009 => x"00000016", --padding
				10010 => x"00000016", --padding
				10011 => x"00000016", --padding
				10012 => x"00000016", --padding
				10013 => x"00000016", --padding
				10014 => x"00000016", --padding
				10015 => x"00000016", --padding
				10016 => x"00000016", --padding
				10017 => x"00000016", --padding
				10018 => x"00000016", --padding
				10019 => x"00000016", --padding
				10020 => x"00000016", --padding
				10021 => x"00000016", --padding
				10022 => x"00000016", --padding
				10023 => x"00000016", --padding
				10024 => x"00000016", --padding
				10025 => x"00000016", --padding
				10026 => x"00000016", --padding
				10027 => x"00000016", --padding
				10028 => x"00000016", --padding
				10029 => x"00000016", --padding
				10030 => x"00000016", --padding
				10031 => x"00000016", --padding
				10032 => x"00000016", --padding
				10033 => x"00000016", --padding
				10034 => x"00000016", --padding
				10035 => x"00000016", --padding
				10036 => x"00000016", --padding
				10037 => x"00000016", --padding
				10038 => x"00000016", --padding
				10039 => x"00000016", --padding
				10040 => x"00000016", --padding
				10041 => x"00000016", --padding
				10042 => x"00000016", --padding
				10043 => x"00000016", --padding
				10044 => x"00000016", --padding
				10045 => x"00000016", --padding
				10046 => x"00000016", --padding
				10047 => x"00000016", --padding
				10048 => x"00000016", --padding
				10049 => x"00000016", --padding
				10050 => x"00000016", --padding
				10051 => x"00000016", --padding
				10052 => x"00000016", --padding
				10053 => x"00000016", --padding
				10054 => x"00000016", --padding
				10055 => x"00000016", --padding
				10056 => x"00000016", --padding
				10057 => x"00000016", --padding
				10058 => x"00000016", --padding
				10059 => x"00000016", --padding
				10060 => x"00000016", --padding
				10061 => x"00000016", --padding
				10062 => x"00000016", --padding
				10063 => x"00000016", --padding
				10064 => x"00000016", --padding
				10065 => x"00000016", --padding
				10066 => x"00000016", --padding
				10067 => x"00000016", --padding
				10068 => x"00000016", --padding
				10069 => x"00000016", --padding
				10070 => x"00000016", --padding
				10071 => x"00000016", --padding
				10072 => x"00000016", --padding
				10073 => x"00000016", --padding
				10074 => x"00000016", --padding
				10075 => x"00000016", --padding
				10076 => x"00000016", --padding
				10077 => x"00000016", --padding
				10078 => x"00000016", --padding
				10079 => x"00000016", --padding
				10080 => x"00000016", --padding
				10081 => x"00000016", --padding
				10082 => x"00000016", --padding
				10083 => x"00000016", --padding
				10084 => x"00000016", --padding
				10085 => x"00000016", --padding
				10086 => x"00000016", --padding
				10087 => x"00000016", --padding
				10088 => x"00000016", --padding
				10089 => x"00000016", --padding
				10090 => x"00000016", --padding
				10091 => x"00000016", --padding
				10092 => x"00000016", --padding
				10093 => x"00000016", --padding
				10094 => x"00000016", --padding
				10095 => x"00000016", --padding
				10096 => x"00000016", --padding
				10097 => x"00000016", --padding
				10098 => x"00000016", --padding
				10099 => x"00000016", --padding
				10100 => x"00000016", --padding
				10101 => x"00000016", --padding
				10102 => x"00000016", --padding
				10103 => x"00000016", --padding
				10104 => x"00000016", --padding
				10105 => x"00000016", --padding
				10106 => x"00000016", --padding
				10107 => x"00000016", --padding
				10108 => x"00000016", --padding
				10109 => x"00000016", --padding
				10110 => x"00000016", --padding
				10111 => x"00000016", --padding
				10112 => x"00000016", --padding
				10113 => x"00000016", --padding
				10114 => x"00000016", --padding
				10115 => x"00000016", --padding
				10116 => x"00000016", --padding
				10117 => x"00000016", --padding
				10118 => x"00000016", --padding
				10119 => x"00000016", --padding
				10120 => x"00000016", --padding
				10121 => x"00000016", --padding
				10122 => x"00000016", --padding
				10123 => x"00000016", --padding
				10124 => x"00000016", --padding
				10125 => x"00000016", --padding
				10126 => x"00000016", --padding
				10127 => x"00000016", --padding
				10128 => x"00000016", --padding
				10129 => x"00000016", --padding
				10130 => x"00000016", --padding
				10131 => x"00000016", --padding
				10132 => x"00000016", --padding
				10133 => x"00000016", --padding
				10134 => x"00000016", --padding
				10135 => x"00000016", --padding
				10136 => x"00000016", --padding
				10137 => x"00000016", --padding
				10138 => x"00000016", --padding
				10139 => x"00000016", --padding
				10140 => x"00000016", --padding
				10141 => x"00000016", --padding
				10142 => x"00000016", --padding
				10143 => x"00000016", --padding
				10144 => x"00000016", --padding
				10145 => x"00000016", --padding
				10146 => x"00000016", --padding
				10147 => x"00000016", --padding
				10148 => x"00000016", --padding
				10149 => x"00000016", --padding
				10150 => x"00000016", --padding
				10151 => x"00000016", --padding
				10152 => x"00000016", --padding
				10153 => x"00000016", --padding
				10154 => x"00000016", --padding
				10155 => x"00000016", --padding
				10156 => x"00000016", --padding
				10157 => x"00000016", --padding
				10158 => x"00000016", --padding
				10159 => x"00000016", --padding
				10160 => x"00000016", --padding
				10161 => x"00000016", --padding
				10162 => x"00000016", --padding
				10163 => x"00000016", --padding
				10164 => x"00000016", --padding
				10165 => x"00000016", --padding
				10166 => x"00000016", --padding
				10167 => x"00000016", --padding
				10168 => x"00000016", --padding
				10169 => x"00000016", --padding
				10170 => x"00000016", --padding
				10171 => x"00000016", --padding
				10172 => x"00000016", --padding
				10173 => x"00000016", --padding
				10174 => x"00000016", --padding
				10175 => x"00000016", --padding
				10176 => x"00000016", --padding
				10177 => x"00000016", --padding
				10178 => x"00000016", --padding
				10179 => x"00000016", --padding
				10180 => x"00000016", --padding
				10181 => x"00000016", --padding
				10182 => x"00000016", --padding
				10183 => x"00000016", --padding
				10184 => x"00000016", --padding
				10185 => x"00000016", --padding
				10186 => x"00000016", --padding
				10187 => x"00000016", --padding
				10188 => x"00000016", --padding
				10189 => x"00000016", --padding
				10190 => x"00000016", --padding
				10191 => x"00000016", --padding
				10192 => x"00000016", --padding
				10193 => x"00000016", --padding
				10194 => x"00000016", --padding
				10195 => x"00000016", --padding
				10196 => x"00000016", --padding
				10197 => x"00000016", --padding
				10198 => x"00000016", --padding
				10199 => x"00000016", --padding
				10200 => x"00000016", --padding
				10201 => x"00000016", --padding
				10202 => x"00000016", --padding
				10203 => x"00000016", --padding
				10204 => x"00000016", --padding
				10205 => x"00000016", --padding
				10206 => x"00000016", --padding
				10207 => x"00000016", --padding
				10208 => x"00000016", --padding
				10209 => x"00000016", --padding
				10210 => x"00000016", --padding
				10211 => x"00000016", --padding
				10212 => x"00000016", --padding
				10213 => x"00000016", --padding
				10214 => x"00000016", --padding
				10215 => x"00000016", --padding
				10216 => x"00000016", --padding
				10217 => x"00000016", --padding
				10218 => x"00000016", --padding
				10219 => x"00000016", --padding
				10220 => x"00000016", --padding
				10221 => x"00000016", --padding
				10222 => x"00000016", --padding
				10223 => x"00000016", --padding
				10224 => x"00000016", --padding
				10225 => x"00000016", --padding
				10226 => x"00000016", --padding
				10227 => x"00000016", --padding
				10228 => x"00000016", --padding
				10229 => x"00000016", --padding
				10230 => x"00000016", --padding
				10231 => x"00000016", --padding
				10232 => x"00000016", --padding
				10233 => x"00000016", --padding
				10234 => x"00000016", --padding
				10235 => x"00000016", --padding
				10236 => x"00000016", --padding
				10237 => x"00000016", --padding
				10238 => x"00000016", --padding
				10239 => x"00000016", --padding
				10240 => x"00000016", --padding
				10241 => x"00000016", --padding
				10242 => x"00000016", --padding
				10243 => x"00000016", --padding
				10244 => x"00000016", --padding
				10245 => x"00000016", --padding
				10246 => x"00000016", --padding
				10247 => x"00000016", --padding
				10248 => x"00000016", --padding
				10249 => x"00000016", --padding
				10250 => x"00000016", --padding
				10251 => x"00000016", --padding
				10252 => x"00000016", --padding
				10253 => x"00000016", --padding
				10254 => x"00000016", --padding
				10255 => x"00000016", --padding
				10256 => x"00000016", --padding
				10257 => x"00000016", --padding
				10258 => x"00000016", --padding
				10259 => x"00000016", --padding
				10260 => x"00000016", --padding
				10261 => x"00000016", --padding
				10262 => x"00000016", --padding
				10263 => x"00000016", --padding
				10264 => x"00000016", --padding
				10265 => x"00000016", --padding
				10266 => x"00000016", --padding
				10267 => x"00000016", --padding
				10268 => x"00000016", --padding
				10269 => x"00000016", --padding
				10270 => x"00000016", --padding
				10271 => x"00000016", --padding
				10272 => x"00000016", --padding
				10273 => x"00000016", --padding
				10274 => x"00000016", --padding
				10275 => x"00000016", --padding
				10276 => x"00000016", --padding
				10277 => x"00000016", --padding
				10278 => x"00000016", --padding
				10279 => x"00000016", --padding
				10280 => x"00000016", --padding
				10281 => x"00000016", --padding
				10282 => x"00000016", --padding
				10283 => x"00000016", --padding
				10284 => x"00000016", --padding
				10285 => x"00000016", --padding
				10286 => x"00000016", --padding
				10287 => x"00000016", --padding
				10288 => x"00000016", --padding
				10289 => x"00000016", --padding
				10290 => x"00000016", --padding
				10291 => x"00000016", --padding
				10292 => x"00000016", --padding
				10293 => x"00000016", --padding
				10294 => x"00000016", --padding
				10295 => x"00000016", --padding
				10296 => x"00000016", --padding
				10297 => x"00000016", --padding
				10298 => x"00000016", --padding
				10299 => x"00000016", --padding
				10300 => x"00000016", --padding
				10301 => x"00000016", --padding
				10302 => x"00000016", --padding
				10303 => x"00000016", --padding
				10304 => x"00000016", --padding
				10305 => x"00000016", --padding
				10306 => x"00000016", --padding
				10307 => x"00000016", --padding
				10308 => x"00000016", --padding
				10309 => x"00000016", --padding
				10310 => x"00000016", --padding
				10311 => x"00000016", --padding
				10312 => x"00000016", --padding
				10313 => x"00000016", --padding
				10314 => x"00000016", --padding
				10315 => x"00000016", --padding
				10316 => x"00000016", --padding
				10317 => x"00000016", --padding
				10318 => x"00000016", --padding
				10319 => x"00000016", --padding
				10320 => x"00000016", --padding
				10321 => x"00000016", --padding
				10322 => x"00000016", --padding
				10323 => x"00000016", --padding
				10324 => x"00000016", --padding
				10325 => x"00000016", --padding
				10326 => x"00000016", --padding
				10327 => x"00000016", --padding
				10328 => x"00000016", --padding
				10329 => x"00000016", --padding
				10330 => x"00000016", --padding
				10331 => x"00000016", --padding
				10332 => x"00000016", --padding
				10333 => x"00000016", --padding
				10334 => x"00000016", --padding
				10335 => x"00000016", --padding
				10336 => x"00000016", --padding
				10337 => x"00000016", --padding
				10338 => x"00000016", --padding
				10339 => x"00000016", --padding
				10340 => x"00000016", --padding
				10341 => x"00000016", --padding
				10342 => x"00000016", --padding
				10343 => x"00000016", --padding
				10344 => x"00000016", --padding
				10345 => x"00000016", --padding
				10346 => x"00000016", --padding
				10347 => x"00000016", --padding
				10348 => x"00000016", --padding
				10349 => x"00000016", --padding
				10350 => x"00000016", --padding
				10351 => x"00000016", --padding
				10352 => x"00000016", --padding
				10353 => x"00000016", --padding
				10354 => x"00000016", --padding
				10355 => x"00000016", --padding
				10356 => x"00000016", --padding
				10357 => x"00000016", --padding
				10358 => x"00000016", --padding
				10359 => x"00000016", --padding
				10360 => x"00000016", --padding
				10361 => x"00000016", --padding
				10362 => x"00000016", --padding
				10363 => x"00000016", --padding
				10364 => x"00000016", --padding
				10365 => x"00000016", --padding
				10366 => x"00000016", --padding
				10367 => x"00000016", --padding
				10368 => x"00000016", --padding
				10369 => x"00000016", --padding
				10370 => x"00000016", --padding
				10371 => x"00000016", --padding
				10372 => x"00000016", --padding
				10373 => x"00000016", --padding
				10374 => x"00000016", --padding
				10375 => x"00000016", --padding
				10376 => x"00000016", --padding
				10377 => x"00000016", --padding
				10378 => x"00000016", --padding
				10379 => x"00000016", --padding
				10380 => x"00000016", --padding
				10381 => x"00000016", --padding
				10382 => x"00000016", --padding
				10383 => x"00000016", --padding
				10384 => x"00000016", --padding
				10385 => x"00000016", --padding
				10386 => x"00000016", --padding
				10387 => x"00000016", --padding
				10388 => x"00000016", --padding
				10389 => x"00000016", --padding
				10390 => x"00000016", --padding
				10391 => x"00000016", --padding
				10392 => x"00000016", --padding
				10393 => x"00000016", --padding
				10394 => x"00000016", --padding
				10395 => x"00000016", --padding
				10396 => x"00000016", --padding
				10397 => x"00000016", --padding
				10398 => x"00000016", --padding
				10399 => x"00000016", --padding
				10400 => x"00000016", --padding
				10401 => x"00000016", --padding
				10402 => x"00000016", --padding
				10403 => x"00000016", --padding
				10404 => x"00000016", --padding
				10405 => x"00000016", --padding
				10406 => x"00000016", --padding
				10407 => x"00000016", --padding
				10408 => x"00000016", --padding
				10409 => x"00000016", --padding
				10410 => x"00000016", --padding
				10411 => x"00000016", --padding
				10412 => x"00000016", --padding
				10413 => x"00000016", --padding
				10414 => x"00000016", --padding
				10415 => x"00000016", --padding
				10416 => x"00000016", --padding
				10417 => x"00000016", --padding
				10418 => x"00000016", --padding
				10419 => x"00000016", --padding
				10420 => x"00000016", --padding
				10421 => x"00000016", --padding
				10422 => x"00000016", --padding
				10423 => x"00000016", --padding
				10424 => x"00000016", --padding
				10425 => x"00000016", --padding
				10426 => x"00000016", --padding
				10427 => x"00000016", --padding
				10428 => x"00000016", --padding
				10429 => x"00000016", --padding
				10430 => x"00000016", --padding
				10431 => x"00000016", --padding
				10432 => x"00000016", --padding
				10433 => x"00000016", --padding
				10434 => x"00000016", --padding
				10435 => x"00000016", --padding
				10436 => x"00000016", --padding
				10437 => x"00000016", --padding
				10438 => x"00000016", --padding
				10439 => x"00000016", --padding
				10440 => x"00000016", --padding
				10441 => x"00000016", --padding
				10442 => x"00000016", --padding
				10443 => x"00000016", --padding
				10444 => x"00000016", --padding
				10445 => x"00000016", --padding
				10446 => x"00000016", --padding
				10447 => x"00000016", --padding
				10448 => x"00000016", --padding
				10449 => x"00000016", --padding
				10450 => x"00000016", --padding
				10451 => x"00000016", --padding
				10452 => x"00000016", --padding
				10453 => x"00000016", --padding
				10454 => x"00000016", --padding
				10455 => x"00000016", --padding
				10456 => x"00000016", --padding
				10457 => x"00000016", --padding
				10458 => x"00000016", --padding
				10459 => x"00000016", --padding
				10460 => x"00000016", --padding
				10461 => x"00000016", --padding
				10462 => x"00000016", --padding
				10463 => x"00000016", --padding
				10464 => x"00000016", --padding
				10465 => x"00000016", --padding
				10466 => x"00000016", --padding
				10467 => x"00000016", --padding
				10468 => x"00000016", --padding
				10469 => x"00000016", --padding
				10470 => x"00000016", --padding
				10471 => x"00000016", --padding
				10472 => x"00000016", --padding
				10473 => x"00000016", --padding
				10474 => x"00000016", --padding
				10475 => x"00000016", --padding
				10476 => x"00000016", --padding
				10477 => x"00000016", --padding
				10478 => x"00000016", --padding
				10479 => x"00000016", --padding
				10480 => x"00000016", --padding
				10481 => x"00000016", --padding
				10482 => x"00000016", --padding
				10483 => x"00000016", --padding
				10484 => x"00000016", --padding
				10485 => x"00000016", --padding
				10486 => x"00000016", --padding
				10487 => x"00000016", --padding
				10488 => x"00000016", --padding
				10489 => x"00000016", --padding
				10490 => x"00000016", --padding
				10491 => x"00000016", --padding
				10492 => x"00000016", --padding
				10493 => x"00000016", --padding
				10494 => x"00000016", --padding
				10495 => x"00000016", --padding
				10496 => x"00000016", --padding
				10497 => x"00000016", --padding
				10498 => x"00000016", --padding
				10499 => x"00000016", --padding
				10500 => x"00000016", --padding
				10501 => x"00000016", --padding
				10502 => x"00000016", --padding
				10503 => x"00000016", --padding
				10504 => x"00000016", --padding
				10505 => x"00000016", --padding
				10506 => x"00000016", --padding
				10507 => x"00000016", --padding
				10508 => x"00000016", --padding
				10509 => x"00000016", --padding
				10510 => x"00000016", --padding
				10511 => x"00000016", --padding
				10512 => x"00000016", --padding
				10513 => x"00000016", --padding
				10514 => x"00000016", --padding
				10515 => x"00000016", --padding
				10516 => x"00000016", --padding
				10517 => x"00000016", --padding
				10518 => x"00000016", --padding
				10519 => x"00000016", --padding
				10520 => x"00000016", --padding
				10521 => x"00000016", --padding
				10522 => x"00000016", --padding
				10523 => x"00000016", --padding
				10524 => x"00000016", --padding
				10525 => x"00000016", --padding
				10526 => x"00000016", --padding
				10527 => x"00000016", --padding
				10528 => x"00000016", --padding
				10529 => x"00000016", --padding
				10530 => x"00000016", --padding
				10531 => x"00000016", --padding
				10532 => x"00000016", --padding
				10533 => x"00000016", --padding
				10534 => x"00000016", --padding
				10535 => x"00000016", --padding
				10536 => x"00000016", --padding
				10537 => x"00000016", --padding
				10538 => x"00000016", --padding
				10539 => x"00000016", --padding
				10540 => x"00000016", --padding
				10541 => x"00000016", --padding
				10542 => x"00000016", --padding
				10543 => x"00000016", --padding
				10544 => x"00000016", --padding
				10545 => x"00000016", --padding
				10546 => x"00000016", --padding
				10547 => x"00000016", --padding
				10548 => x"00000016", --padding
				10549 => x"00000016", --padding
				10550 => x"00000016", --padding
				10551 => x"00000016", --padding
				10552 => x"00000016", --padding
				10553 => x"00000016", --padding
				10554 => x"00000016", --padding
				10555 => x"00000016", --padding
				10556 => x"00000016", --padding
				10557 => x"00000016", --padding
				10558 => x"00000016", --padding
				10559 => x"00000016", --padding
				10560 => x"00000016", --padding
				10561 => x"00000016", --padding
				10562 => x"00000016", --padding
				10563 => x"00000016", --padding
				10564 => x"00000016", --padding
				10565 => x"00000016", --padding
				10566 => x"00000016", --padding
				10567 => x"00000016", --padding
				10568 => x"00000016", --padding
				10569 => x"00000016", --padding
				10570 => x"00000016", --padding
				10571 => x"00000016", --padding
				10572 => x"00000016", --padding
				10573 => x"00000016", --padding
				10574 => x"00000016", --padding
				10575 => x"00000016", --padding
				10576 => x"00000016", --padding
				10577 => x"00000016", --padding
				10578 => x"00000016", --padding
				10579 => x"00000016", --padding
				10580 => x"00000016", --padding
				10581 => x"00000016", --padding
				10582 => x"00000016", --padding
				10583 => x"00000016", --padding
				10584 => x"00000016", --padding
				10585 => x"00000016", --padding
				10586 => x"00000016", --padding
				10587 => x"00000016", --padding
				10588 => x"00000016", --padding
				10589 => x"00000016", --padding
				10590 => x"00000016", --padding
				10591 => x"00000016", --padding
				10592 => x"00000016", --padding
				10593 => x"00000016", --padding
				10594 => x"00000016", --padding
				10595 => x"00000016", --padding
				10596 => x"00000016", --padding
				10597 => x"00000016", --padding
				10598 => x"00000016", --padding
				10599 => x"00000016", --padding
				10600 => x"00000016", --padding
				10601 => x"00000016", --padding
				10602 => x"00000016", --padding
				10603 => x"00000016", --padding
				10604 => x"00000016", --padding
				10605 => x"00000016", --padding
				10606 => x"00000016", --padding
				10607 => x"00000016", --padding
				10608 => x"00000016", --padding
				10609 => x"00000016", --padding
				10610 => x"00000016", --padding
				10611 => x"00000016", --padding
				10612 => x"00000016", --padding
				10613 => x"00000016", --padding
				10614 => x"00000016", --padding
				10615 => x"00000016", --padding
				10616 => x"00000016", --padding
				10617 => x"00000016", --padding
				10618 => x"00000016", --padding
				10619 => x"00000016", --padding
				10620 => x"00000016", --padding
				10621 => x"00000016", --padding
				10622 => x"00000016", --padding
				10623 => x"00000016", --padding
				10624 => x"00000016", --padding
				10625 => x"00000016", --padding
				10626 => x"00000016", --padding
				10627 => x"00000016", --padding
				10628 => x"00000016", --padding
				10629 => x"00000016", --padding
				10630 => x"00000016", --padding
				10631 => x"00000016", --padding
				10632 => x"00000016", --padding
				10633 => x"00000016", --padding
				10634 => x"00000016", --padding
				10635 => x"00000016", --padding
				10636 => x"00000016", --padding
				10637 => x"00000016", --padding
				10638 => x"00000016", --padding
				10639 => x"00000016", --padding
				10640 => x"00000016", --padding
				10641 => x"00000016", --padding
				10642 => x"00000016", --padding
				10643 => x"00000016", --padding
				10644 => x"00000016", --padding
				10645 => x"00000016", --padding
				10646 => x"00000016", --padding
				10647 => x"00000016", --padding
				10648 => x"00000016", --padding
				10649 => x"00000016", --padding
				10650 => x"00000016", --padding
				10651 => x"00000016", --padding
				10652 => x"00000016", --padding
				10653 => x"00000016", --padding
				10654 => x"00000016", --padding
				10655 => x"00000016", --padding
				10656 => x"00000016", --padding
				10657 => x"00000016", --padding
				10658 => x"00000016", --padding
				10659 => x"00000016", --padding
				10660 => x"00000016", --padding
				10661 => x"00000016", --padding
				10662 => x"00000016", --padding
				10663 => x"00000016", --padding
				10664 => x"00000016", --padding
				10665 => x"00000016", --padding
				10666 => x"00000016", --padding
				10667 => x"00000016", --padding
				10668 => x"00000016", --padding
				10669 => x"00000016", --padding
				10670 => x"00000016", --padding
				10671 => x"00000016", --padding
				10672 => x"00000016", --padding
				10673 => x"00000016", --padding
				10674 => x"00000016", --padding
				10675 => x"00000016", --padding
				10676 => x"00000016", --padding
				10677 => x"00000016", --padding
				10678 => x"00000016", --padding
				10679 => x"00000016", --padding
				10680 => x"00000016", --padding
				10681 => x"00000016", --padding
				10682 => x"00000016", --padding
				10683 => x"00000016", --padding
				10684 => x"00000016", --padding
				10685 => x"00000016", --padding
				10686 => x"00000016", --padding
				10687 => x"00000016", --padding
				10688 => x"00000016", --padding
				10689 => x"00000016", --padding
				10690 => x"00000016", --padding
				10691 => x"00000016", --padding
				10692 => x"00000016", --padding
				10693 => x"00000016", --padding
				10694 => x"00000016", --padding
				10695 => x"00000016", --padding
				10696 => x"00000016", --padding
				10697 => x"00000016", --padding
				10698 => x"00000016", --padding
				10699 => x"00000016", --padding
				10700 => x"00000016", --padding
				10701 => x"00000016", --padding
				10702 => x"00000016", --padding
				10703 => x"00000016", --padding
				10704 => x"00000016", --padding
				10705 => x"00000016", --padding
				10706 => x"00000016", --padding
				10707 => x"00000016", --padding
				10708 => x"00000016", --padding
				10709 => x"00000016", --padding
				10710 => x"00000016", --padding
				10711 => x"00000016", --padding
				10712 => x"00000016", --padding
				10713 => x"00000016", --padding
				10714 => x"00000016", --padding
				10715 => x"00000016", --padding
				10716 => x"00000016", --padding
				10717 => x"00000016", --padding
				10718 => x"00000016", --padding
				10719 => x"00000016", --padding
				10720 => x"00000016", --padding
				10721 => x"00000016", --padding
				10722 => x"00000016", --padding
				10723 => x"00000016", --padding
				10724 => x"00000016", --padding
				10725 => x"00000016", --padding
				10726 => x"00000016", --padding
				10727 => x"00000016", --padding
				10728 => x"00000016", --padding
				10729 => x"00000016", --padding
				10730 => x"00000016", --padding
				10731 => x"00000016", --padding
				10732 => x"00000016", --padding
				10733 => x"00000016", --padding
				10734 => x"00000016", --padding
				10735 => x"00000016", --padding
				10736 => x"00000016", --padding
				10737 => x"00000016", --padding
				10738 => x"00000016", --padding
				10739 => x"00000016", --padding
				10740 => x"00000016", --padding
				10741 => x"00000016", --padding
				10742 => x"00000016", --padding
				10743 => x"00000016", --padding
				10744 => x"00000016", --padding
				10745 => x"00000016", --padding
				10746 => x"00000016", --padding
				10747 => x"00000016", --padding
				10748 => x"00000016", --padding
				10749 => x"00000016", --padding
				10750 => x"00000016", --padding
				10751 => x"00000016", --padding
				10752 => x"00000016", --padding
				10753 => x"00000016", --padding
				10754 => x"00000016", --padding
				10755 => x"00000016", --padding
				10756 => x"00000016", --padding
				10757 => x"00000016", --padding
				10758 => x"00000016", --padding
				10759 => x"00000016", --padding
				10760 => x"00000016", --padding
				10761 => x"00000016", --padding
				10762 => x"00000016", --padding
				10763 => x"00000016", --padding
				10764 => x"00000016", --padding
				10765 => x"00000016", --padding
				10766 => x"00000016", --padding
				10767 => x"00000016", --padding
				10768 => x"00000016", --padding
				10769 => x"00000016", --padding
				10770 => x"00000016", --padding
				10771 => x"00000016", --padding
				10772 => x"00000016", --padding
				10773 => x"00000016", --padding
				10774 => x"00000016", --padding
				10775 => x"00000016", --padding
				10776 => x"00000016", --padding
				10777 => x"00000016", --padding
				10778 => x"00000016", --padding
				10779 => x"00000016", --padding
				10780 => x"00000016", --padding
				10781 => x"00000016", --padding
				10782 => x"00000016", --padding
				10783 => x"00000016", --padding
				10784 => x"00000016", --padding
				10785 => x"00000016", --padding
				10786 => x"00000016", --padding
				10787 => x"00000016", --padding
				10788 => x"00000016", --padding
				10789 => x"00000016", --padding
				10790 => x"00000016", --padding
				10791 => x"00000016", --padding
				10792 => x"00000016", --padding
				10793 => x"00000016", --padding
				10794 => x"00000016", --padding
				10795 => x"00000016", --padding
				10796 => x"00000016", --padding
				10797 => x"00000016", --padding
				10798 => x"00000016", --padding
				10799 => x"00000016", --padding
				10800 => x"00000016", --padding
				10801 => x"00000016", --padding
				10802 => x"00000016", --padding
				10803 => x"00000016", --padding
				10804 => x"00000016", --padding
				10805 => x"00000016", --padding
				10806 => x"00000016", --padding
				10807 => x"00000016", --padding
				10808 => x"00000016", --padding
				10809 => x"00000016", --padding
				10810 => x"00000016", --padding
				10811 => x"00000016", --padding
				10812 => x"00000016", --padding
				10813 => x"00000016", --padding
				10814 => x"00000016", --padding
				10815 => x"00000016", --padding
				10816 => x"00000016", --padding
				10817 => x"00000016", --padding
				10818 => x"00000016", --padding
				10819 => x"00000016", --padding
				10820 => x"00000016", --padding
				10821 => x"00000016", --padding
				10822 => x"00000016", --padding
				10823 => x"00000016", --padding
				10824 => x"00000016", --padding
				10825 => x"00000016", --padding
				10826 => x"00000016", --padding
				10827 => x"00000016", --padding
				10828 => x"00000016", --padding
				10829 => x"00000016", --padding
				10830 => x"00000016", --padding
				10831 => x"00000016", --padding
				10832 => x"00000016", --padding
				10833 => x"00000016", --padding
				10834 => x"00000016", --padding
				10835 => x"00000016", --padding
				10836 => x"00000016", --padding
				10837 => x"00000016", --padding
				10838 => x"00000016", --padding
				10839 => x"00000016", --padding
				10840 => x"00000016", --padding
				10841 => x"00000016", --padding
				10842 => x"00000016", --padding
				10843 => x"00000016", --padding
				10844 => x"00000016", --padding
				10845 => x"00000016", --padding
				10846 => x"00000016", --padding
				10847 => x"00000016", --padding
				10848 => x"00000016", --padding
				10849 => x"00000016", --padding
				10850 => x"00000016", --padding
				10851 => x"00000016", --padding
				10852 => x"00000016", --padding
				10853 => x"00000016", --padding
				10854 => x"00000016", --padding
				10855 => x"00000016", --padding
				10856 => x"00000016", --padding
				10857 => x"00000016", --padding
				10858 => x"00000016", --padding
				10859 => x"00000016", --padding
				10860 => x"00000016", --padding
				10861 => x"00000016", --padding
				10862 => x"00000016", --padding
				10863 => x"00000016", --padding
				10864 => x"00000016", --padding
				10865 => x"00000016", --padding
				10866 => x"00000016", --padding
				10867 => x"00000016", --padding
				10868 => x"00000016", --padding
				10869 => x"00000016", --padding
				10870 => x"00000016", --padding
				10871 => x"00000016", --padding
				10872 => x"00000016", --padding
				10873 => x"00000016", --padding
				10874 => x"00000016", --padding
				10875 => x"00000016", --padding
				10876 => x"00000016", --padding
				10877 => x"00000016", --padding
				10878 => x"00000016", --padding
				10879 => x"00000016", --padding
				10880 => x"00000016", --padding
				10881 => x"00000016", --padding
				10882 => x"00000016", --padding
				10883 => x"00000016", --padding
				10884 => x"00000016", --padding
				10885 => x"00000016", --padding
				10886 => x"00000016", --padding
				10887 => x"00000016", --padding
				10888 => x"00000016", --padding
				10889 => x"00000016", --padding
				10890 => x"00000016", --padding
				10891 => x"00000016", --padding
				10892 => x"00000016", --padding
				10893 => x"00000016", --padding
				10894 => x"00000016", --padding
				10895 => x"00000016", --padding
				10896 => x"00000016", --padding
				10897 => x"00000016", --padding
				10898 => x"00000016", --padding
				10899 => x"00000016", --padding
				10900 => x"00000016", --padding
				10901 => x"00000016", --padding
				10902 => x"00000016", --padding
				10903 => x"00000016", --padding
				10904 => x"00000016", --padding
				10905 => x"00000016", --padding
				10906 => x"00000016", --padding
				10907 => x"00000016", --padding
				10908 => x"00000016", --padding
				10909 => x"00000016", --padding
				10910 => x"00000016", --padding
				10911 => x"00000016", --padding
				10912 => x"00000016", --padding
				10913 => x"00000016", --padding
				10914 => x"00000016", --padding
				10915 => x"00000016", --padding
				10916 => x"00000016", --padding
				10917 => x"00000016", --padding
				10918 => x"00000016", --padding
				10919 => x"00000016", --padding
				10920 => x"00000016", --padding
				10921 => x"00000016", --padding
				10922 => x"00000016", --padding
				10923 => x"00000016", --padding
				10924 => x"00000016", --padding
				10925 => x"00000016", --padding
				10926 => x"00000016", --padding
				10927 => x"00000016", --padding
				10928 => x"00000016", --padding
				10929 => x"00000016", --padding
				10930 => x"00000016", --padding
				10931 => x"00000016", --padding
				10932 => x"00000016", --padding
				10933 => x"00000016", --padding
				10934 => x"00000016", --padding
				10935 => x"00000016", --padding
				10936 => x"00000016", --padding
				10937 => x"00000016", --padding
				10938 => x"00000016", --padding
				10939 => x"00000016", --padding
				10940 => x"00000016", --padding
				10941 => x"00000016", --padding
				10942 => x"00000016", --padding
				10943 => x"00000016", --padding
				10944 => x"00000016", --padding
				10945 => x"00000016", --padding
				10946 => x"00000016", --padding
				10947 => x"00000016", --padding
				10948 => x"00000016", --padding
				10949 => x"00000016", --padding
				10950 => x"00000016", --padding
				10951 => x"00000016", --padding
				10952 => x"00000016", --padding
				10953 => x"00000016", --padding
				10954 => x"00000016", --padding
				10955 => x"00000016", --padding
				10956 => x"00000016", --padding
				10957 => x"00000016", --padding
				10958 => x"00000016", --padding
				10959 => x"00000016", --padding
				10960 => x"00000016", --padding
				10961 => x"00000016", --padding
				10962 => x"00000016", --padding
				10963 => x"00000016", --padding
				10964 => x"00000016", --padding
				10965 => x"00000016", --padding
				10966 => x"00000016", --padding
				10967 => x"00000016", --padding
				10968 => x"00000016", --padding
				10969 => x"00000016", --padding
				10970 => x"00000016", --padding
				10971 => x"00000016", --padding
				10972 => x"00000016", --padding
				10973 => x"00000016", --padding
				10974 => x"00000016", --padding
				10975 => x"00000016", --padding
				10976 => x"00000016", --padding
				10977 => x"00000016", --padding
				10978 => x"00000016", --padding
				10979 => x"00000016", --padding
				10980 => x"00000016", --padding
				10981 => x"00000016", --padding
				10982 => x"00000016", --padding
				10983 => x"00000016", --padding
				10984 => x"00000016", --padding
				10985 => x"00000016", --padding
				10986 => x"00000016", --padding
				10987 => x"00000016", --padding
				10988 => x"00000016", --padding
				10989 => x"00000016", --padding
				10990 => x"00000016", --padding
				10991 => x"00000016", --padding
				10992 => x"00000016", --padding
				10993 => x"00000016", --padding
				10994 => x"00000016", --padding
				10995 => x"00000016", --padding
				10996 => x"00000016", --padding
				10997 => x"00000016", --padding
				10998 => x"00000016", --padding
				10999 => x"00000016", --padding
				11000 => x"00000016", --padding
				11001 => x"00000016", --padding
				11002 => x"00000016", --padding
				11003 => x"00000016", --padding
				11004 => x"00000016", --padding
				11005 => x"00000016", --padding
				11006 => x"00000016", --padding
				11007 => x"00000016", --padding
				11008 => x"00000016", --padding
				11009 => x"00000016", --padding
				11010 => x"00000016", --padding
				11011 => x"00000016", --padding
				11012 => x"00000016", --padding
				11013 => x"00000016", --padding
				11014 => x"00000016", --padding
				11015 => x"00000016", --padding
				11016 => x"00000016", --padding
				11017 => x"00000016", --padding
				11018 => x"00000016", --padding
				11019 => x"00000016", --padding
				11020 => x"00000016", --padding
				11021 => x"00000016", --padding
				11022 => x"00000016", --padding
				11023 => x"00000016", --padding
				11024 => x"00000016", --padding
				11025 => x"00000016", --padding
				11026 => x"00000016", --padding
				11027 => x"00000016", --padding
				11028 => x"00000016", --padding
				11029 => x"00000016", --padding
				11030 => x"00000016", --padding
				11031 => x"00000016", --padding
				11032 => x"00000016", --padding
				11033 => x"00000016", --padding
				11034 => x"00000016", --padding
				11035 => x"00000016", --padding
				11036 => x"00000016", --padding
				11037 => x"00000016", --padding
				11038 => x"00000016", --padding
				11039 => x"00000016", --padding
				11040 => x"00000016", --padding
				11041 => x"00000016", --padding
				11042 => x"00000016", --padding
				11043 => x"00000016", --padding
				11044 => x"00000016", --padding
				11045 => x"00000016", --padding
				11046 => x"00000016", --padding
				11047 => x"00000016", --padding
				11048 => x"00000016", --padding
				11049 => x"00000016", --padding
				11050 => x"00000016", --padding
				11051 => x"00000016", --padding
				11052 => x"00000016", --padding
				11053 => x"00000016", --padding
				11054 => x"00000016", --padding
				11055 => x"00000016", --padding
				11056 => x"00000016", --padding
				11057 => x"00000016", --padding
				11058 => x"00000016", --padding
				11059 => x"00000016", --padding
				11060 => x"00000016", --padding
				11061 => x"00000016", --padding
				11062 => x"00000016", --padding
				11063 => x"00000016", --padding
				11064 => x"00000016", --padding
				11065 => x"00000016", --padding
				11066 => x"00000016", --padding
				11067 => x"00000016", --padding
				11068 => x"00000016", --padding
				11069 => x"00000016", --padding
				11070 => x"00000016", --padding
				11071 => x"00000016", --padding
				11072 => x"00000016", --padding
				11073 => x"00000016", --padding
				11074 => x"00000016", --padding
				11075 => x"00000016", --padding
				11076 => x"00000016", --padding
				11077 => x"00000016", --padding
				11078 => x"00000016", --padding
				11079 => x"00000016", --padding
				11080 => x"00000016", --padding
				11081 => x"00000016", --padding
				11082 => x"00000016", --padding
				11083 => x"00000016", --padding
				11084 => x"00000016", --padding
				11085 => x"00000016", --padding
				11086 => x"00000016", --padding
				11087 => x"00000016", --padding
				11088 => x"00000016", --padding
				11089 => x"00000016", --padding
				11090 => x"00000016", --padding
				11091 => x"00000016", --padding
				11092 => x"00000016", --padding
				11093 => x"00000016", --padding
				11094 => x"00000016", --padding
				11095 => x"00000016", --padding
				11096 => x"00000016", --padding
				11097 => x"00000016", --padding
				11098 => x"00000016", --padding
				11099 => x"00000016", --padding
				11100 => x"00000016", --padding
				11101 => x"00000016", --padding
				11102 => x"00000016", --padding
				11103 => x"00000016", --padding
				11104 => x"00000016", --padding
				11105 => x"00000016", --padding
				11106 => x"00000016", --padding
				11107 => x"00000016", --padding
				11108 => x"00000016", --padding
				11109 => x"00000016", --padding
				11110 => x"00000016", --padding
				11111 => x"00000016", --padding
				11112 => x"00000016", --padding
				11113 => x"00000016", --padding
				11114 => x"00000016", --padding
				11115 => x"00000016", --padding
				11116 => x"00000016", --padding
				11117 => x"00000016", --padding
				11118 => x"00000016", --padding
				11119 => x"00000016", --padding
				11120 => x"00000016", --padding
				11121 => x"00000016", --padding
				11122 => x"00000016", --padding
				11123 => x"00000016", --padding
				11124 => x"00000016", --padding
				11125 => x"00000016", --padding
				11126 => x"00000016", --padding
				11127 => x"00000016", --padding
				11128 => x"00000016", --padding
				11129 => x"00000016", --padding
				11130 => x"00000016", --padding
				11131 => x"00000016", --padding
				11132 => x"00000016", --padding
				11133 => x"00000016", --padding
				11134 => x"00000016", --padding
				11135 => x"00000016", --padding
				11136 => x"00000016", --padding
				11137 => x"00000016", --padding
				11138 => x"00000016", --padding
				11139 => x"00000016", --padding
				11140 => x"00000016", --padding
				11141 => x"00000016", --padding
				11142 => x"00000016", --padding
				11143 => x"00000016", --padding
				11144 => x"00000016", --padding
				11145 => x"00000016", --padding
				11146 => x"00000016", --padding
				11147 => x"00000016", --padding
				11148 => x"00000016", --padding
				11149 => x"00000016", --padding
				11150 => x"00000016", --padding
				11151 => x"00000016", --padding
				11152 => x"00000016", --padding
				11153 => x"00000016", --padding
				11154 => x"00000016", --padding
				11155 => x"00000016", --padding
				11156 => x"00000016", --padding
				11157 => x"00000016", --padding
				11158 => x"00000016", --padding
				11159 => x"00000016", --padding
				11160 => x"00000016", --padding
				11161 => x"00000016", --padding
				11162 => x"00000016", --padding
				11163 => x"00000016", --padding
				11164 => x"00000016", --padding
				11165 => x"00000016", --padding
				11166 => x"00000016", --padding
				11167 => x"00000016", --padding
				11168 => x"00000016", --padding
				11169 => x"00000016", --padding
				11170 => x"00000016", --padding
				11171 => x"00000016", --padding
				11172 => x"00000016", --padding
				11173 => x"00000016", --padding
				11174 => x"00000016", --padding
				11175 => x"00000016", --padding
				11176 => x"00000016", --padding
				11177 => x"00000016", --padding
				11178 => x"00000016", --padding
				11179 => x"00000016", --padding
				11180 => x"00000016", --padding
				11181 => x"00000016", --padding
				11182 => x"00000016", --padding

				----------------------------------------------------

others => x"00000000"
	);


begin

	process(i_clk)
	begin
		if rising_edge(i_clk) then
			-- memory write --
			if i_we = '1' then
				mem(to_integer(unsigned(i_w_addr))) <= i_data;
			end if;
			-- memory read --
			o_data <= mem(to_integer(unsigned(i_r_addr)));

		end if;
	end process;

end architecture arch;
